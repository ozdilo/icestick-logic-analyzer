-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2016.02.27810

-- Build Date:         Jan 29 2016 01:59:39

-- File Generated:     Aug 24 2016 00:01:56

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "la" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of la
entity la is
port (
    debugleds : out std_logic_vector(1 downto 0);
    testcnt : out std_logic_vector(7 downto 0);
    input : in std_logic_vector(7 downto 0);
    xtalClock : in std_logic;
    tx : out std_logic;
    rx : in std_logic;
    ready50 : out std_logic;
    exClock : in std_logic);
end la;

-- Architecture of la
-- View name is \INTERFACE\
architecture \INTERFACE\ of la is

signal \N__38006\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \VCCG0\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_6\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_5\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_4\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_3\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_2\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_7\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_8\ : std_logic;
signal \n234_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_9\ : std_logic;
signal n234 : std_logic;
signal \byteDone\ : std_logic;
signal \n9_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.bits_3\ : std_logic;
signal \Inst_eia232.Inst_transmitter.bits_2\ : std_logic;
signal n3493 : std_logic;
signal \n3493_cascade_\ : std_logic;
signal n6749 : std_logic;
signal \Inst_eia232.Inst_transmitter.bits_0\ : std_logic;
signal \Inst_eia232.Inst_transmitter.bits_1\ : std_logic;
signal n4082 : std_logic;
signal \Inst_eia232.Inst_transmitter.counter_3\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n2201_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.counter_4\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n8642\ : std_logic;
signal \Inst_eia232.Inst_transmitter.counter_1\ : std_logic;
signal \Inst_eia232.Inst_transmitter.counter_2\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n3594\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n3594_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n4719\ : std_logic;
signal n3615 : std_logic;
signal \Inst_eia232.Inst_transmitter.counter_0\ : std_logic;
signal outputdata_0 : std_logic;
signal outputdata_4 : std_logic;
signal outputdata_5 : std_logic;
signal \Inst_eia232.Inst_transmitter.txBuffer_1\ : std_logic;
signal tx_c : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7836\ : std_logic;
signal \GENERIC_FIFO_1.n7837\ : std_logic;
signal \GENERIC_FIFO_1.n7838\ : std_logic;
signal \GENERIC_FIFO_1.n7839\ : std_logic;
signal \GENERIC_FIFO_1.n7840\ : std_logic;
signal \GENERIC_FIFO_1.n7841\ : std_logic;
signal \GENERIC_FIFO_1.n7842\ : std_logic;
signal \GENERIC_FIFO_1.n7843\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7844\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7827\ : std_logic;
signal \GENERIC_FIFO_1.n7828\ : std_logic;
signal \GENERIC_FIFO_1.n7829\ : std_logic;
signal \GENERIC_FIFO_1.n7830\ : std_logic;
signal \GENERIC_FIFO_1.n7831\ : std_logic;
signal \GENERIC_FIFO_1.n7832\ : std_logic;
signal \GENERIC_FIFO_1.n7833\ : std_logic;
signal \GENERIC_FIFO_1.n7834\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7835\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_7\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_1\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_4\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_3\ : std_logic;
signal \GENERIC_FIFO_1.n12\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \GENERIC_FIFO_1.n11\ : std_logic;
signal \GENERIC_FIFO_1.n7818\ : std_logic;
signal \GENERIC_FIFO_1.n10\ : std_logic;
signal \GENERIC_FIFO_1.n7819\ : std_logic;
signal \GENERIC_FIFO_1.n9\ : std_logic;
signal \GENERIC_FIFO_1.n7820\ : std_logic;
signal \GENERIC_FIFO_1.n8\ : std_logic;
signal \GENERIC_FIFO_1.n7821\ : std_logic;
signal \GENERIC_FIFO_1.n7\ : std_logic;
signal \GENERIC_FIFO_1.n7822\ : std_logic;
signal \GENERIC_FIFO_1.n6\ : std_logic;
signal \GENERIC_FIFO_1.n7823\ : std_logic;
signal \GENERIC_FIFO_1.n5\ : std_logic;
signal \GENERIC_FIFO_1.n7824\ : std_logic;
signal \GENERIC_FIFO_1.n7825\ : std_logic;
signal \GENERIC_FIFO_1.n4\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7826\ : std_logic;
signal \GENERIC_FIFO_1.n3\ : std_logic;
signal \n4005_cascade_\ : std_logic;
signal \dataBuffer_22\ : std_logic;
signal \dataBuffer_30\ : std_logic;
signal \dataBuffer_24\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_0\ : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_8\ : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_0\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n3571\ : std_logic;
signal \dataBuffer_19\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n8854_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_3\ : std_logic;
signal \dataBuffer_14\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n1323\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n3632_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_6\ : std_logic;
signal \dataBuffer_18\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n8851_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_2\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_1\ : std_logic;
signal \n4248_cascade_\ : std_logic;
signal \n1336_cascade_\ : std_logic;
signal \dataBuffer_25\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n8847\ : std_logic;
signal n4248 : std_logic;
signal n1320 : std_logic;
signal \n1320_cascade_\ : std_logic;
signal \dataBuffer_28\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n8756_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_4\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_4\ : std_logic;
signal \state_1_N_371_1_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n1\ : std_logic;
signal bytes_1 : std_logic;
signal bytes_2 : std_logic;
signal \Inst_eia232.Inst_transmitter.n9218_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n3\ : std_logic;
signal disabled : std_logic;
signal \Inst_eia232.Inst_transmitter.n6745\ : std_logic;
signal \state_1_N_371_1\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n3652\ : std_logic;
signal bytes_0 : std_logic;
signal \Inst_eia232.Inst_transmitter.n3652_cascade_\ : std_logic;
signal n1336 : std_logic;
signal outputdata_1 : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_1\ : std_logic;
signal outputdata_2 : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_2\ : std_logic;
signal outputdata_3 : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_3\ : std_logic;
signal outputdata_6 : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_6\ : std_logic;
signal \Inst_eia232.Inst_transmitter.disabledBuffer_1\ : std_logic;
signal \disabledGroupsReg_1\ : std_logic;
signal \Inst_eia232.Inst_transmitter.disabledBuffer_3\ : std_logic;
signal \disabledGroupsReg_3\ : std_logic;
signal \Inst_eia232.Inst_transmitter.disabledBuffer_2\ : std_logic;
signal \disabledGroupsReg_2\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_7\ : std_logic;
signal outputdata_7 : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_7\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7929\ : std_logic;
signal \GENERIC_FIFO_1.n7930\ : std_logic;
signal \GENERIC_FIFO_1.n7931\ : std_logic;
signal \GENERIC_FIFO_1.n7932\ : std_logic;
signal \GENERIC_FIFO_1.n7933\ : std_logic;
signal \GENERIC_FIFO_1.n7934\ : std_logic;
signal \GENERIC_FIFO_1.n7935\ : std_logic;
signal \GENERIC_FIFO_1.n7936\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7937\ : std_logic;
signal \maskRegister_5\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n6703\ : std_logic;
signal \Inst_eia232.Inst_transmitter.dataBuffer_5\ : std_logic;
signal \Inst_eia232.Inst_transmitter.byte_5\ : std_logic;
signal \GENERIC_FIFO_1.n8677_cascade_\ : std_logic;
signal \GENERIC_FIFO_1.n1396_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4743\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_0\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_8\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_9\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_7\ : std_logic;
signal \GENERIC_FIFO_1.n18_cascade_\ : std_logic;
signal \GENERIC_FIFO_1.fifo_memory_N_983\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n11\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_5\ : std_logic;
signal \GENERIC_FIFO_1.n16_cascade_\ : std_logic;
signal \GENERIC_FIFO_1.n20_adj_1274\ : std_logic;
signal \GENERIC_FIFO_1.n4721\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_925_0\ : std_logic;
signal \GENERIC_FIFO_1.n24\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \GENERIC_FIFO_1.n23\ : std_logic;
signal \GENERIC_FIFO_1.n7809\ : std_logic;
signal \GENERIC_FIFO_1.n22\ : std_logic;
signal \GENERIC_FIFO_1.n7810\ : std_logic;
signal \GENERIC_FIFO_1.n21\ : std_logic;
signal \GENERIC_FIFO_1.n7811\ : std_logic;
signal \GENERIC_FIFO_1.n20\ : std_logic;
signal \GENERIC_FIFO_1.n7812\ : std_logic;
signal \GENERIC_FIFO_1.n19\ : std_logic;
signal \GENERIC_FIFO_1.n7813\ : std_logic;
signal \GENERIC_FIFO_1.n18_adj_1275\ : std_logic;
signal \GENERIC_FIFO_1.n7814\ : std_logic;
signal \GENERIC_FIFO_1.n17\ : std_logic;
signal \GENERIC_FIFO_1.n7815\ : std_logic;
signal \GENERIC_FIFO_1.n7816\ : std_logic;
signal \GENERIC_FIFO_1.n16_adj_1273\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \GENERIC_FIFO_1.n7817\ : std_logic;
signal \GENERIC_FIFO_1.n15\ : std_logic;
signal \GENERIC_FIFO_1.n8650\ : std_logic;
signal \GENERIC_FIFO_1.n8681\ : std_logic;
signal \GENERIC_FIFO_1.n78\ : std_logic;
signal \GENERIC_FIFO_1.level_9__N_900\ : std_logic;
signal \GENERIC_FIFO_1.n8654\ : std_logic;
signal \GENERIC_FIFO_1.n1418\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_6\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_2\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_6\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_0\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_8\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_5\ : std_logic;
signal \GENERIC_FIFO_1.n16_adj_1276_cascade_\ : std_logic;
signal \GENERIC_FIFO_1.level_9_N_876_9\ : std_logic;
signal \GENERIC_FIFO_1.n17_adj_1278\ : std_logic;
signal \GENERIC_FIFO_1.n1396\ : std_logic;
signal \GENERIC_FIFO_1.n18_adj_1277\ : std_logic;
signal \GENERIC_FIFO_1.n141_cascade_\ : std_logic;
signal \GENERIC_FIFO_1.n69\ : std_logic;
signal \Inst_eia232.Inst_receiver.n2143_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.bitcount_1\ : std_logic;
signal \Inst_eia232.Inst_receiver.bitcount_2\ : std_logic;
signal \Inst_eia232.Inst_receiver.bitcount_3\ : std_logic;
signal \Inst_eia232.Inst_receiver.bitcount_0\ : std_logic;
signal \Inst_eia232.Inst_receiver.n7_adj_1264_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8769_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n6736_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8772\ : std_logic;
signal \Inst_eia232.Inst_receiver.bytecount_2\ : std_logic;
signal \Inst_eia232.Inst_receiver.bytecount_1\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8582_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8831_cascade_\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n3552\ : std_logic;
signal \Inst_eia232.xon\ : std_logic;
signal \Inst_eia232.Inst_receiver.n75_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n5597\ : std_logic;
signal \Inst_eia232.Inst_receiver.n5597_cascade_\ : std_logic;
signal \Inst_eia232.xoff\ : std_logic;
signal \Inst_eia232.Inst_receiver.n90_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n5498\ : std_logic;
signal cmd_6 : std_logic;
signal \n5698_cascade_\ : std_logic;
signal \nstate_2_N_241_0\ : std_logic;
signal \Inst_eia232.Inst_receiver.n14_adj_1265\ : std_logic;
signal \Inst_eia232.Inst_receiver.n112\ : std_logic;
signal \Inst_eia232.Inst_receiver.n112_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n90\ : std_logic;
signal \GENERIC_FIFO_1.n8779\ : std_logic;
signal \valueRegister_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n9114_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n9108\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6\ : std_logic;
signal \GENERIC_FIFO_1.n71\ : std_logic;
signal \GENERIC_FIFO_1.n70\ : std_logic;
signal \Inst_eia232.Inst_receiver.n4628\ : std_logic;
signal \Inst_eia232.Inst_transmitter.paused\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n4634\ : std_logic;
signal state_0 : std_logic;
signal \Inst_eia232.Inst_transmitter.n2580\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n8527\ : std_logic;
signal \Inst_eia232.id\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n971\ : std_logic;
signal state_1 : std_logic;
signal \Inst_eia232.Inst_transmitter.n4712\ : std_logic;
signal \GENERIC_FIFO_1.n77\ : std_logic;
signal \GENERIC_FIFO_1.n76\ : std_logic;
signal \GENERIC_FIFO_1.n75\ : std_logic;
signal \GENERIC_FIFO_1.n74\ : std_logic;
signal \GENERIC_FIFO_1.n73\ : std_logic;
signal \GENERIC_FIFO_1.n1420\ : std_logic;
signal \GENERIC_FIFO_1.n72\ : std_logic;
signal \GENERIC_FIFO_1.n16_adj_1279_cascade_\ : std_logic;
signal \GENERIC_FIFO_1.n142\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_7\ : std_logic;
signal \GENERIC_FIFO_1.n17_adj_1280\ : std_logic;
signal \GENERIC_FIFO_1.n1421\ : std_logic;
signal \GENERIC_FIFO_1.n1423\ : std_logic;
signal \writeByte\ : std_logic;
signal n9 : std_logic;
signal \Inst_eia232.Inst_transmitter.n3608\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_0\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_1\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_2\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_3\ : std_logic;
signal \GENERIC_FIFO_1.write_pointer_6\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_0\ : std_logic;
signal \GENERIC_FIFO_1.n2\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \GENERIC_FIFO_1.n1379\ : std_logic;
signal \GENERIC_FIFO_1.n7938\ : std_logic;
signal \GENERIC_FIFO_1.n1391\ : std_logic;
signal \GENERIC_FIFO_1.n1378\ : std_logic;
signal \GENERIC_FIFO_1.n8634\ : std_logic;
signal \GENERIC_FIFO_1.n7939\ : std_logic;
signal \GENERIC_FIFO_1.n1377\ : std_logic;
signal \GENERIC_FIFO_1.n7940\ : std_logic;
signal \GENERIC_FIFO_1.n1390\ : std_logic;
signal \GENERIC_FIFO_1.n1376\ : std_logic;
signal \GENERIC_FIFO_1.n8628\ : std_logic;
signal \GENERIC_FIFO_1.n7941\ : std_logic;
signal \GENERIC_FIFO_1.n1375\ : std_logic;
signal \GENERIC_FIFO_1.n7942\ : std_logic;
signal \GENERIC_FIFO_1.n1386\ : std_logic;
signal \GENERIC_FIFO_1.n1374\ : std_logic;
signal \GENERIC_FIFO_1.n8632\ : std_logic;
signal \GENERIC_FIFO_1.n7943\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \GENERIC_FIFO_1.n7944\ : std_logic;
signal \GENERIC_FIFO_1.n7944_THRU_CRY_0_THRU_CO\ : std_logic;
signal \GENERIC_FIFO_1.n1388\ : std_logic;
signal \GENERIC_FIFO_1.n1373\ : std_logic;
signal \GENERIC_FIFO_1.n8630\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \GENERIC_FIFO_1.n1372\ : std_logic;
signal \GENERIC_FIFO_1.n7945\ : std_logic;
signal \GENERIC_FIFO_1.n1383\ : std_logic;
signal \GENERIC_FIFO_1.n1371\ : std_logic;
signal \GENERIC_FIFO_1.n8638\ : std_logic;
signal \GENERIC_FIFO_1.n7946\ : std_logic;
signal \GENERIC_FIFO_1.n1392\ : std_logic;
signal \GENERIC_FIFO_1.n1392_THRU_CO\ : std_logic;
signal \GENERIC_FIFO_1.n8821\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_9\ : std_logic;
signal \GENERIC_FIFO_1.n1416\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8755_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n9123_cascade_\ : std_logic;
signal \executePrev\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8784\ : std_logic;
signal \Inst_eia232.Inst_receiver.n6_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n5504\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8782_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n6_adj_1267\ : std_logic;
signal \Inst_eia232.Inst_receiver.n3_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n5505\ : std_logic;
signal \Inst_eia232.Inst_receiver.n3504_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.n3676\ : std_logic;
signal \Inst_eia232.Inst_receiver.n4767\ : std_logic;
signal \Inst_eia232.Inst_receiver.n3504\ : std_logic;
signal \Inst_eia232.Inst_receiver.n5\ : std_logic;
signal \Inst_eia232.Inst_receiver.n75\ : std_logic;
signal \Inst_eia232.Inst_receiver.n14\ : std_logic;
signal n1917 : std_logic;
signal \Inst_eia232.Inst_receiver.counter_4\ : std_logic;
signal \Inst_eia232.Inst_receiver.counter_3\ : std_logic;
signal \Inst_eia232.Inst_receiver.n7_cascade_\ : std_logic;
signal \Inst_eia232.Inst_receiver.counter_1\ : std_logic;
signal \Inst_eia232.Inst_receiver.counter_0\ : std_logic;
signal \Inst_eia232.Inst_receiver.counter_2\ : std_logic;
signal \Inst_eia232.Inst_receiver.n7777\ : std_logic;
signal \Inst_eia232.Inst_receiver.n3202\ : std_logic;
signal \Inst_eia232.Inst_receiver.n1_adj_1266\ : std_logic;
signal \Inst_eia232.state_0\ : std_logic;
signal \Inst_eia232.Inst_receiver.nstate_2_N_133_1\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8826\ : std_logic;
signal \Inst_eia232.Inst_prescaler.counter_4__N_38\ : std_logic;
signal \Inst_eia232.Inst_receiver.cmd_4\ : std_logic;
signal \Inst_eia232.Inst_receiver.cmd_5\ : std_logic;
signal n12 : std_logic;
signal \Inst_eia232.Inst_receiver.cmd_1\ : std_logic;
signal \Inst_eia232.Inst_receiver.n3718\ : std_logic;
signal \Inst_eia232.Inst_receiver.cmd_2\ : std_logic;
signal \Inst_eia232.Inst_receiver.cmd_0\ : std_logic;
signal \Inst_eia232.Inst_receiver.cmd_3\ : std_logic;
signal \Inst_eia232.Inst_receiver.n69\ : std_logic;
signal \Inst_eia232.state_1\ : std_logic;
signal \Inst_eia232.state_2\ : std_logic;
signal \Inst_eia232.Inst_prescaler.counter_1\ : std_logic;
signal \Inst_eia232.Inst_prescaler.counter_0\ : std_logic;
signal \trxClock\ : std_logic;
signal \nstate_2__N_139_c_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n9096_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_cascade_\ : std_logic;
signal \configRegister_23_adj_1379\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n9102_cascade_\ : std_logic;
signal \valueRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n9084_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_cascade_\ : std_logic;
signal \configRegister_23_adj_1339\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n9090_cascade_\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4730\ : std_logic;
signal \valueRegister_2\ : std_logic;
signal \valueRegister_5\ : std_logic;
signal \configRegister_24\ : std_logic;
signal \maskRegister_0_adj_1288\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4642\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_1\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_2\ : std_logic;
signal \valueRegister_6\ : std_logic;
signal \maskRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4740\ : std_logic;
signal \maskRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4741\ : std_logic;
signal \maskRegister_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4742\ : std_logic;
signal \maskRegister_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4744\ : std_logic;
signal \maskRegister_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4745\ : std_logic;
signal \valueRegister_4\ : std_logic;
signal \GENERIC_FIFO_1.n1422\ : std_logic;
signal \valueRegister_7\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4729\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_4\ : std_logic;
signal \GENERIC_FIFO_1.n8815\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_3\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4731\ : std_logic;
signal \GENERIC_FIFO_1.n1424\ : std_logic;
signal \GENERIC_FIFO_1.n1419\ : std_logic;
signal \GENERIC_FIFO_1.n8813\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_1\ : std_logic;
signal \GENERIC_FIFO_1.n8814\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_2\ : std_logic;
signal \GENERIC_FIFO_1.n1417\ : std_logic;
signal \GENERIC_FIFO_1.n8816\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_4\ : std_logic;
signal \GENERIC_FIFO_1.n8817\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_5\ : std_logic;
signal \GENERIC_FIFO_1.n8818\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_6\ : std_logic;
signal \GENERIC_FIFO_1.n8819\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_7\ : std_logic;
signal \GENERIC_FIFO_1.n141\ : std_logic;
signal \GENERIC_FIFO_1.n8820\ : std_logic;
signal \GENERIC_FIFO_1.read_pointer_8\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_0\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4732\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input180Delay_4\ : std_logic;
signal testcnt_c_0 : std_logic;
signal \bfn_6_1_0_\ : std_logic;
signal testcnt_c_1 : std_logic;
signal n7862 : std_logic;
signal testcnt_c_2 : std_logic;
signal n7863 : std_logic;
signal testcnt_c_3 : std_logic;
signal n7864 : std_logic;
signal testcnt_c_4 : std_logic;
signal n7865 : std_logic;
signal testcnt_c_5 : std_logic;
signal n7866 : std_logic;
signal testcnt_c_6 : std_logic;
signal n7867 : std_logic;
signal n7868 : std_logic;
signal testcnt_c_7 : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \configRegister_1_adj_1399\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7914\ : std_logic;
signal \configRegister_2_adj_1398\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7915\ : std_logic;
signal \configRegister_3_adj_1397\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7916\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7917\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7918\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7919\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7920\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7921\ : std_logic;
signal \configRegister_8_adj_1392\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7922\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7923\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7924\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7925\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7926\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7927\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7928\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15\ : std_logic;
signal \Inst_eia232.Inst_receiver.n7_adj_1264\ : std_logic;
signal \Inst_eia232.Inst_receiver.n957\ : std_logic;
signal \Inst_eia232.Inst_receiver.bytecount_0\ : std_logic;
signal \Inst_eia232.Inst_receiver.n3557\ : std_logic;
signal \Inst_eia232.Inst_receiver.n8376\ : std_logic;
signal \maskRegister_6_adj_1362\ : std_logic;
signal \maskRegister_7_adj_1361\ : std_logic;
signal \maskRegister_4_adj_1364\ : std_logic;
signal \configRegister_6_adj_1394\ : std_logic;
signal \maskRegister_3_adj_1365\ : std_logic;
signal \configRegister_7_adj_1393\ : std_logic;
signal \valueRegister_0_adj_1296\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_3\ : std_logic;
signal \configRegister_0_adj_1400\ : std_logic;
signal \configRegister_20_adj_1342\ : std_logic;
signal \configRegister_4_adj_1396\ : std_logic;
signal cmd_39 : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4641\ : std_logic;
signal \configRegister_21_adj_1381\ : std_logic;
signal wrtrigval_0 : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1\ : std_logic;
signal \valueRegister_1\ : std_logic;
signal \configRegister_26\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n9078\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_cascade_\ : std_logic;
signal \configRegister_21_adj_1301\ : std_logic;
signal \configRegister_23_adj_1299\ : std_logic;
signal \configRegister_22_adj_1300\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n9072_cascade_\ : std_logic;
signal \configRegister_20_adj_1302\ : std_logic;
signal \configRegister_24_adj_1298\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0\ : std_logic;
signal \maskRegister_1_adj_1287\ : std_logic;
signal \maskRegister_2_adj_1286\ : std_logic;
signal \maskRegister_3_adj_1285\ : std_logic;
signal \maskRegister_5_adj_1283\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_2\ : std_logic;
signal \Inst_core.Inst_sync.n2789_cascade_\ : std_logic;
signal \syncedInput_2\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_6\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_6\ : std_logic;
signal \maskRegister_4_adj_1284\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4637\ : std_logic;
signal \maskRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4739\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input180Delay_7\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_5\ : std_logic;
signal \Inst_core.Inst_sync.n9063_cascade_\ : std_logic;
signal \syncedInput_5\ : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput_4\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_4\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_4\ : std_logic;
signal \Inst_core.Inst_sync.n9057_cascade_\ : std_logic;
signal \syncedInput_4\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input180Delay_6\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4734\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input180Delay_5\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4733\ : std_logic;
signal input_c_4 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_4\ : std_logic;
signal \INVInst_core.Inst_sync.synchronizedInput180_i4C_net\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4765\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n25_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n27\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n26\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4766\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n28\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n28\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n25_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n27\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n26\ : std_logic;
signal \valueRegister_6_adj_1370\ : std_logic;
signal \configRegister_5_adj_1395\ : std_logic;
signal \valueRegister_7_adj_1369\ : std_logic;
signal \configRegister_11_adj_1389\ : std_logic;
signal \configRegister_10_adj_1390\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_7\ : std_logic;
signal \configRegister_15_adj_1385\ : std_logic;
signal \configRegister_24_adj_1378\ : std_logic;
signal \Inst_eia232.Inst_transmitter.n4246\ : std_logic;
signal n4005 : std_logic;
signal \disabledGroupsReg_0\ : std_logic;
signal \Inst_eia232.Inst_transmitter.disabledBuffer_0\ : std_logic;
signal \configRegister_22_adj_1380\ : std_logic;
signal \configRegister_23\ : std_logic;
signal wrtrigmask_0 : std_logic;
signal \maskRegister_0\ : std_logic;
signal \configRegister_20_adj_1382\ : std_logic;
signal \configRegister_22_adj_1340\ : std_logic;
signal \configRegister_21\ : std_logic;
signal wrtrigmask_1 : std_logic;
signal \configRegister_21_adj_1341\ : std_logic;
signal \wrFlags\ : std_logic;
signal cmd_32 : std_logic;
signal \configRegister_20\ : std_logic;
signal \valueRegister_1_adj_1295\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4746\ : std_logic;
signal fwd_15 : std_logic;
signal \Inst_core.Inst_controller.n22_cascade_\ : std_logic;
signal fwd_6 : std_logic;
signal \Inst_core.Inst_controller.n4_adj_986_cascade_\ : std_logic;
signal fwd_5 : std_logic;
signal \Inst_core.Inst_controller.n4_adj_987_cascade_\ : std_logic;
signal \Inst_core.Inst_controller.n8486\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_0\ : std_logic;
signal \syncedInput_3\ : std_logic;
signal \syncedInput_7\ : std_logic;
signal \valueRegister_7_adj_1329\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_1\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_3\ : std_logic;
signal \Inst_core.Inst_sync.n2791\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_0\ : std_logic;
signal \Inst_core.Inst_sync.n2793\ : std_logic;
signal \flagInverted\ : std_logic;
signal \flagFilter\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_1\ : std_logic;
signal \Inst_core.Inst_sync.n2787\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_5\ : std_logic;
signal \syncedInput_6\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_6\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_7\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_2\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_5\ : std_logic;
signal \Inst_core.Inst_sync.n9117\ : std_logic;
signal \Inst_core.Inst_sync.demuxedInput_3\ : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput_5\ : std_logic;
signal \Inst_core.Inst_sync.n2566\ : std_logic;
signal \Inst_core.Inst_sync.n2564\ : std_logic;
signal \Inst_core.Inst_sync.n9129\ : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput_6\ : std_logic;
signal input_c_0 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_0\ : std_logic;
signal input_c_1 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_1\ : std_logic;
signal input_c_2 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_2\ : std_logic;
signal input_c_3 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_3\ : std_logic;
signal input_c_6 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_6\ : std_logic;
signal input_c_5 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_5\ : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput180_7\ : std_logic;
signal \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\ : std_logic;
signal \Inst_core.n8518_cascade_\ : std_logic;
signal \valueRegister_7_adj_1289\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_7\ : std_logic;
signal \memoryOut_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n8808_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n3\ : std_logic;
signal \Inst_core.n1639_cascade_\ : std_logic;
signal \Inst_core.n9054\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \configRegister_1_adj_1359\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7899\ : std_logic;
signal \configRegister_2_adj_1358\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7900\ : std_logic;
signal \configRegister_3_adj_1357\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7901\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7902\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7903\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7904\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7905\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7906\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7907\ : std_logic;
signal \configRegister_10_adj_1350\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7908\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7909\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7910\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7911\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7912\ : std_logic;
signal \Inst_core.n1639\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7913\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4114\ : std_logic;
signal \Inst_core.configRegister_27\ : std_logic;
signal \configRegister_7_adj_1353\ : std_logic;
signal \configRegister_11_adj_1349\ : std_logic;
signal \configRegister_12_adj_1388\ : std_logic;
signal \configRegister_5_adj_1355\ : std_logic;
signal \configRegister_14_adj_1346\ : std_logic;
signal \configRegister_9_adj_1351\ : std_logic;
signal \configRegister_8_adj_1352\ : std_logic;
signal cmd_16 : std_logic;
signal \configRegister_15_adj_1345\ : std_logic;
signal wrtrigmask_3 : std_logic;
signal \configRegister_9_adj_1391\ : std_logic;
signal cmd_38 : std_logic;
signal \Inst_core.Inst_controller.fwd_14\ : std_logic;
signal cmd_30 : std_logic;
signal \configRegister_22\ : std_logic;
signal cmd_33 : std_logic;
signal cmd_37 : std_logic;
signal cmd_36 : std_logic;
signal \configRegister_6_adj_1354\ : std_logic;
signal \valueRegister_5_adj_1291\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4750\ : std_logic;
signal bwd_11 : std_logic;
signal bwd_8 : std_logic;
signal fwd_11 : std_logic;
signal fwd_4 : std_logic;
signal \Inst_core.Inst_controller.n18_cascade_\ : std_logic;
signal \Inst_core.Inst_controller.n21\ : std_logic;
signal fwd_13 : std_logic;
signal fwd_9 : std_logic;
signal \Inst_core.Inst_controller.n15\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4\ : std_logic;
signal \valueRegister_4_adj_1292\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4749\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_4\ : std_logic;
signal fwd_12 : std_logic;
signal fwd_1 : std_logic;
signal \Inst_core.Inst_controller.n13\ : std_logic;
signal bwd_10 : std_logic;
signal \Inst_core.Inst_controller.n14\ : std_logic;
signal fwd_8 : std_logic;
signal \Inst_core.Inst_controller.n11\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n14\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n11\ : std_logic;
signal cmd_29 : std_logic;
signal \syncedInput_0\ : std_logic;
signal \syncedInput_1\ : std_logic;
signal \valueRegister_4_adj_1332\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4756\ : std_logic;
signal \Inst_core.Inst_sampler.n31_adj_995_cascade_\ : std_logic;
signal divider_9 : std_logic;
signal divider_7 : std_logic;
signal \Inst_core.Inst_sampler.n29\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_4\ : std_logic;
signal \valueRegister_5_adj_1331\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_5\ : std_logic;
signal divider_15 : std_logic;
signal divider_13 : std_logic;
signal divider_16 : std_logic;
signal \Inst_core.Inst_sampler.n32\ : std_logic;
signal divider_14 : std_logic;
signal \Inst_core.Inst_sampler.n8596_cascade_\ : std_logic;
signal \Inst_core.Inst_sampler.n8590\ : std_logic;
signal \valueRegister_1_adj_1335\ : std_logic;
signal divider_20 : std_logic;
signal divider_21 : std_logic;
signal \Inst_core.Inst_sampler.n8598\ : std_logic;
signal \Inst_core.Inst_sampler.n8602\ : std_logic;
signal \Inst_core.Inst_sampler.n8600_cascade_\ : std_logic;
signal \Inst_core.Inst_sampler.n8604\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelL16\ : std_logic;
signal \configRegister_24_adj_1338\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n8844_cascade_\ : std_logic;
signal \Inst_core.Inst_decoder.n6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n9052\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n1765\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n667\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n667_cascade_\ : std_logic;
signal \Inst_core.n31_adj_1174\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n100_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n656\ : std_logic;
signal \Inst_core.n8518\ : std_logic;
signal \Inst_core.state_1_adj_1134\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n657\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n554\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n22_cascade_\ : std_logic;
signal \Inst_core.n8515_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n451\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n760\ : std_logic;
signal \Inst_core.n31\ : std_logic;
signal cmd_18 : std_logic;
signal \configRegister_13_adj_1347\ : std_logic;
signal \configRegister_14_adj_1386\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5\ : std_logic;
signal \memoryOut_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n2_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n100\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n553\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n100_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n2_cascade_\ : std_logic;
signal \configRegister_17_adj_1383\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n100\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n100_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n759\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n770\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.state_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n770_cascade_\ : std_logic;
signal \Inst_core.n6713\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4076\ : std_logic;
signal \configRegister_17_adj_1303\ : std_logic;
signal \configRegister_4_adj_1356\ : std_logic;
signal \maskRegister_5_adj_1363\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4764\ : std_logic;
signal \configRegister_12_adj_1348\ : std_logic;
signal \Inst_core.arm\ : std_logic;
signal \maskRegister_5_adj_1323\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4757\ : std_logic;
signal \maskRegister_6_adj_1322\ : std_logic;
signal \maskRegister_7_adj_1321\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4759\ : std_logic;
signal \maskRegister_0_adj_1368\ : std_logic;
signal \maskRegister_1_adj_1367\ : std_logic;
signal \maskRegister_2_adj_1366\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7_adj_996\ : std_logic;
signal \flagDemux\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register\ : std_logic;
signal \valueRegister_5_adj_1371\ : std_logic;
signal \configRegister_13_adj_1387\ : std_logic;
signal wrtrigcfg_3 : std_logic;
signal \configRegister_16_adj_1384\ : std_logic;
signal \configRegister_16_adj_1304\ : std_logic;
signal cmd_17 : std_logic;
signal cmd_28 : std_logic;
signal fwd_3 : std_logic;
signal bwd_9 : std_logic;
signal \Inst_core.Inst_controller.n24\ : std_logic;
signal \Inst_core.Inst_controller.n22_adj_988_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3\ : std_logic;
signal \valueRegister_3_adj_1293\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4748\ : std_logic;
signal bwd_6 : std_logic;
signal bwd_5 : std_logic;
signal \Inst_core.Inst_controller.n23\ : std_logic;
signal bwd_3 : std_logic;
signal bwd_4 : std_logic;
signal \Inst_core.Inst_controller.n21_adj_989\ : std_logic;
signal cmd_11 : std_logic;
signal cmd_15 : std_logic;
signal bwd_7 : std_logic;
signal fwd_10 : std_logic;
signal wrtrigmask_2 : std_logic;
signal \maskRegister_4_adj_1324\ : std_logic;
signal \Inst_core.Inst_sync.filteredInput_7\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.n4735\ : std_logic;
signal \maskRegister_7_adj_1281\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4752\ : std_logic;
signal \maskRegister_0_adj_1328\ : std_logic;
signal \maskRegister_1_adj_1327\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4753\ : std_logic;
signal \maskRegister_2_adj_1326\ : std_logic;
signal \maskRegister_3_adj_1325\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6\ : std_logic;
signal \valueRegister_6_adj_1330\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4758\ : std_logic;
signal divider_4 : std_logic;
signal \Inst_core.Inst_sampler.n30\ : std_logic;
signal \Inst_core.Inst_sampler.n8592\ : std_logic;
signal divider_2 : std_logic;
signal divider_10 : std_logic;
signal divider_8 : std_logic;
signal divider_17 : std_logic;
signal \Inst_core.Inst_sampler.n8588\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \Inst_core.Inst_sampler.n7948\ : std_logic;
signal \Inst_core.Inst_sampler.n7949\ : std_logic;
signal \Inst_core.Inst_sampler.n7950\ : std_logic;
signal \Inst_core.Inst_sampler.counter_4\ : std_logic;
signal \Inst_core.Inst_sampler.n7951\ : std_logic;
signal \Inst_core.Inst_sampler.n7952\ : std_logic;
signal \Inst_core.Inst_sampler.n7953\ : std_logic;
signal \Inst_core.Inst_sampler.counter_7\ : std_logic;
signal \Inst_core.Inst_sampler.n7954\ : std_logic;
signal \Inst_core.Inst_sampler.n7955\ : std_logic;
signal \Inst_core.Inst_sampler.counter_8\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \Inst_core.Inst_sampler.counter_9\ : std_logic;
signal \Inst_core.Inst_sampler.n7956\ : std_logic;
signal \Inst_core.Inst_sampler.counter_10\ : std_logic;
signal \Inst_core.Inst_sampler.n7957\ : std_logic;
signal \Inst_core.Inst_sampler.n7958\ : std_logic;
signal \Inst_core.Inst_sampler.n7959\ : std_logic;
signal \Inst_core.Inst_sampler.counter_13\ : std_logic;
signal \Inst_core.Inst_sampler.n7960\ : std_logic;
signal \Inst_core.Inst_sampler.counter_14\ : std_logic;
signal \Inst_core.Inst_sampler.n7961\ : std_logic;
signal \Inst_core.Inst_sampler.counter_15\ : std_logic;
signal \Inst_core.Inst_sampler.n7962\ : std_logic;
signal \Inst_core.Inst_sampler.n7963\ : std_logic;
signal \Inst_core.Inst_sampler.counter_16\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \Inst_core.Inst_sampler.counter_17\ : std_logic;
signal \Inst_core.Inst_sampler.n7964\ : std_logic;
signal \Inst_core.Inst_sampler.n7965\ : std_logic;
signal \Inst_core.Inst_sampler.counter_19\ : std_logic;
signal \Inst_core.Inst_sampler.n7966\ : std_logic;
signal \Inst_core.Inst_sampler.counter_20\ : std_logic;
signal \Inst_core.Inst_sampler.n7967\ : std_logic;
signal \Inst_core.Inst_sampler.counter_21\ : std_logic;
signal \Inst_core.Inst_sampler.n7968\ : std_logic;
signal \Inst_core.Inst_sampler.n7969\ : std_logic;
signal \Inst_core.Inst_sampler.n7970\ : std_logic;
signal \Inst_core.Inst_sampler.n1700\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n8622\ : std_logic;
signal cmd_35 : std_logic;
signal \configRegister_0_adj_1360\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4\ : std_logic;
signal \memoryOut_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4763\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n11\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n6675_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n564\ : std_logic;
signal \Inst_core.n8837\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.state_1\ : std_logic;
signal \configRegister_0_adj_1320\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n9055\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \configRegister_1_adj_1319\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7884\ : std_logic;
signal \configRegister_2_adj_1318\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7885\ : std_logic;
signal \configRegister_3_adj_1317\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7886\ : std_logic;
signal \configRegister_4_adj_1316\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7887\ : std_logic;
signal \configRegister_5_adj_1315\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7888\ : std_logic;
signal \configRegister_6_adj_1314\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7889\ : std_logic;
signal \configRegister_7_adj_1313\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7890\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7891\ : std_logic;
signal \configRegister_8_adj_1312\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \configRegister_9_adj_1311\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7892\ : std_logic;
signal \configRegister_10_adj_1310\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7893\ : std_logic;
signal \configRegister_11_adj_1309\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7894\ : std_logic;
signal \configRegister_12_adj_1308\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7895\ : std_logic;
signal \configRegister_13_adj_1307\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7896\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7897\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n1662\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n7898\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4144\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4761\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n2_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n100\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n100_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n450\ : std_logic;
signal \Inst_core.Inst_trigger.levelReg_0\ : std_logic;
signal \configRegister_17_adj_1343\ : std_logic;
signal \Inst_core.Inst_trigger.levelReg_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n99\ : std_logic;
signal \valueRegister_4_adj_1372\ : std_logic;
signal \configRegister_15_adj_1305\ : std_logic;
signal bwd_15 : std_logic;
signal \configRegister_17\ : std_logic;
signal cmd_21 : std_logic;
signal wrtrigcfg_1 : std_logic;
signal \configRegister_14_adj_1306\ : std_logic;
signal cmd_12 : std_logic;
signal fwd_7 : std_logic;
signal \maskRegister_6_adj_1282\ : std_logic;
signal cmd_31 : std_logic;
signal cmd_10 : std_logic;
signal \valueRegister_2_adj_1374\ : std_logic;
signal cmd_25 : std_logic;
signal wrtrigval_2 : std_logic;
signal cmd_22 : std_logic;
signal cmd_26 : std_logic;
signal cmd_27 : std_logic;
signal divider_19 : std_logic;
signal bwd_2 : std_logic;
signal bwd_13 : std_logic;
signal \Inst_core.Inst_controller.n18_adj_990\ : std_logic;
signal \Inst_core.Inst_controller.n20\ : std_logic;
signal \Inst_core.Inst_controller.n17_cascade_\ : std_logic;
signal \Inst_core.Inst_controller.n30\ : std_logic;
signal \Inst_core.Inst_controller.n29_cascade_\ : std_logic;
signal \Inst_core.Inst_controller.n6693\ : std_logic;
signal \Inst_core.Inst_controller.bwd_14\ : std_logic;
signal \Inst_core.Inst_controller.n19\ : std_logic;
signal \valueRegister_2_adj_1294\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4747\ : std_logic;
signal \memoryOut_6\ : std_logic;
signal \configRegister_26_adj_1297\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n4751\ : std_logic;
signal fwd_0 : std_logic;
signal fwd_2 : std_logic;
signal \Inst_core.Inst_controller.n16\ : std_logic;
signal debugleds_c_1 : std_logic;
signal \Inst_core.n4_cascade_\ : std_logic;
signal \Inst_core.Inst_controller.n3907_cascade_\ : std_logic;
signal \memoryOut_2\ : std_logic;
signal \valueRegister_2_adj_1334\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4754\ : std_logic;
signal divider_11 : std_logic;
signal \Inst_core.Inst_sampler.counter_23\ : std_logic;
signal \Inst_core.Inst_sampler.counter_11\ : std_logic;
signal \Inst_core.Inst_sampler.counter_2\ : std_logic;
signal \Inst_core.Inst_sampler.n8606\ : std_logic;
signal \Inst_core.Inst_sampler.n3_cascade_\ : std_logic;
signal divider_23 : std_logic;
signal \Inst_core.Inst_sampler.n8618\ : std_logic;
signal \Inst_core.Inst_sampler.n8656_cascade_\ : std_logic;
signal divider_1 : std_logic;
signal \Inst_core.Inst_sampler.counter_18\ : std_logic;
signal divider_18 : std_logic;
signal \Inst_core.Inst_sampler.counter_1\ : std_logic;
signal \Inst_core.Inst_sampler.n28\ : std_logic;
signal \Inst_core.Inst_sampler.n27_cascade_\ : std_logic;
signal divider_6 : std_logic;
signal \Inst_core.Inst_sampler.counter_3\ : std_logic;
signal divider_3 : std_logic;
signal \Inst_core.Inst_sampler.counter_6\ : std_logic;
signal \Inst_core.Inst_sampler.n26\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3\ : std_logic;
signal \valueRegister_3_adj_1333\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4755\ : std_logic;
signal divider_0 : std_logic;
signal \Inst_core.Inst_sampler.counter_12\ : std_logic;
signal divider_12 : std_logic;
signal \Inst_core.Inst_sampler.counter_0\ : std_logic;
signal \Inst_core.Inst_sampler.n25\ : std_logic;
signal \Inst_core.Inst_sync.Inst_filter.input360_7\ : std_logic;
signal input_c_7 : std_logic;
signal \Inst_core.Inst_sync.synchronizedInput_7\ : std_logic;
signal cmd_13 : std_logic;
signal \Inst_core.Inst_sampler.n35\ : std_logic;
signal \Inst_core.Inst_sampler.n36\ : std_logic;
signal \Inst_core.Inst_sampler.n33\ : std_logic;
signal \wrDivider\ : std_logic;
signal \Inst_core.Inst_sampler.n8669\ : std_logic;
signal \Inst_core.Inst_sampler.n8671\ : std_logic;
signal \Inst_core.Inst_sampler.n8673\ : std_logic;
signal \Inst_core.Inst_sampler.n8687\ : std_logic;
signal \valueRegister_0_adj_1336\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n4643\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_2__Inst_stage.n7\ : std_logic;
signal divider_5 : std_logic;
signal \Inst_core.Inst_sampler.counter_22\ : std_logic;
signal divider_22 : std_logic;
signal \Inst_core.Inst_sampler.counter_5\ : std_logic;
signal \Inst_core.Inst_sampler.n34\ : std_logic;
signal \Inst_core.Inst_sampler.n44\ : std_logic;
signal \Inst_core.Inst_sampler.n43\ : std_logic;
signal \Inst_core.Inst_sampler.n45\ : std_logic;
signal \ready50_N_581\ : std_logic;
signal \Inst_core.configRegister_27_adj_1196\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n8626\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4\ : std_logic;
signal \memoryOut_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4645\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7_adj_1000\ : std_logic;
signal \Inst_core.Inst_trigger.configRegister_27\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n8521_cascade_\ : std_logic;
signal \Inst_core.n3670\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n7\ : std_logic;
signal \Inst_core.Inst_trigger.stageRun_0\ : std_logic;
signal \Inst_core.Inst_trigger.stageRun_3\ : std_logic;
signal \Inst_core.stageRun_2\ : std_logic;
signal \Inst_core.stageRun_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n8753_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n461\ : std_logic;
signal \Inst_core.state_1\ : std_logic;
signal \valueRegister_3_adj_1373\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3\ : std_logic;
signal \memoryOut_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4762\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n28\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n25_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n31\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n27\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8\ : std_logic;
signal \Inst_core.Inst_trigger.stages_1__Inst_stage.n26\ : std_logic;
signal \configRegister_0\ : std_logic;
signal \Inst_core.n9053\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7869\ : std_logic;
signal \configRegister_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7870\ : std_logic;
signal \configRegister_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7871\ : std_logic;
signal \configRegister_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7872\ : std_logic;
signal \configRegister_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7873\ : std_logic;
signal \configRegister_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7874\ : std_logic;
signal \configRegister_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7875\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7876\ : std_logic;
signal \configRegister_8\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \configRegister_9\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7877\ : std_logic;
signal \configRegister_10\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7878\ : std_logic;
signal \configRegister_11\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7879\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7880\ : std_logic;
signal \configRegister_13\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7881\ : std_logic;
signal \configRegister_14\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7882\ : std_logic;
signal \Inst_core.n1705\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n7883\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n4044\ : std_logic;
signal \valueRegister_1_adj_1375\ : std_logic;
signal \memoryOut_1\ : std_logic;
signal \configRegister_26_adj_1377\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_3__Inst_stage.n4760\ : std_logic;
signal \Inst_core.Inst_trigger.stageMatch_2\ : std_logic;
signal \Inst_core.Inst_trigger.stageMatch_3\ : std_logic;
signal \Inst_core.Inst_trigger.stageMatch_1\ : std_logic;
signal \Inst_core.Inst_trigger.stageMatch_0\ : std_logic;
signal \Inst_core.Inst_trigger.levelReg_1__N_590\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n28\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n25_cascade_\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n27\ : std_logic;
signal \Inst_core.n31_adj_1132\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3\ : std_logic;
signal \Inst_core.Inst_trigger.stages_0__Inst_stage.n26\ : std_logic;
signal \configRegister_1\ : std_logic;
signal \configRegister_16\ : std_logic;
signal n3753 : std_logic;
signal n1 : std_logic;
signal cmd_19 : std_logic;
signal wrtrigval_1 : std_logic;
signal cmd_14 : std_logic;
signal \valueRegister_6_adj_1290\ : std_logic;
signal \configRegister_12\ : std_logic;
signal cmd_9 : std_logic;
signal bwd_1 : std_logic;
signal wrtrigcfg_0 : std_logic;
signal cmd_23 : std_logic;
signal \configRegister_15\ : std_logic;
signal cmd_24 : std_logic;
signal \configRegister_16_adj_1344\ : std_logic;
signal wrtrigval_3 : std_logic;
signal \valueRegister_0_adj_1376\ : std_logic;
signal cmd_8 : std_logic;
signal bwd_0 : std_logic;
signal wrtrigcfg_2 : std_logic;
signal cmd_34 : std_logic;
signal \configRegister_26_adj_1337\ : std_logic;
signal wrsize : std_logic;
signal cmd_20 : std_logic;
signal bwd_12 : std_logic;
signal \Inst_core.nstate_1_N_831_0\ : std_logic;
signal \Inst_core.Inst_controller.n321\ : std_logic;
signal \Inst_core.Inst_controller.nstate_1_N_827_1\ : std_logic;
signal \Inst_core.resetCmd\ : std_logic;
signal debugleds_c_0 : std_logic;
signal busy : std_logic;
signal \Inst_core.Inst_controller.nstate_1_N_825_0\ : std_logic;
signal \Inst_core.Inst_controller.n320\ : std_logic;
signal \Inst_core.Inst_controller.nstate_1_N_829_0\ : std_logic;
signal \Inst_core.Inst_controller.n2717\ : std_logic;
signal \sampleReady\ : std_logic;
signal \Inst_core.n318\ : std_logic;
signal \Inst_core.Inst_controller.n2717_cascade_\ : std_logic;
signal send : std_logic;
signal \Inst_core.Inst_controller.n2\ : std_logic;
signal \Inst_core.Inst_controller.counter_0\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \Inst_core.Inst_controller.counter_1\ : std_logic;
signal \Inst_core.Inst_controller.n7845\ : std_logic;
signal \Inst_core.Inst_controller.counter_2\ : std_logic;
signal \Inst_core.Inst_controller.n7846\ : std_logic;
signal \Inst_core.Inst_controller.counter_3\ : std_logic;
signal \Inst_core.Inst_controller.n7847\ : std_logic;
signal \Inst_core.Inst_controller.counter_4\ : std_logic;
signal \Inst_core.Inst_controller.n7848\ : std_logic;
signal \Inst_core.Inst_controller.counter_5\ : std_logic;
signal \Inst_core.Inst_controller.n7849\ : std_logic;
signal \Inst_core.Inst_controller.counter_6\ : std_logic;
signal \Inst_core.Inst_controller.n7850\ : std_logic;
signal \Inst_core.Inst_controller.counter_7\ : std_logic;
signal \Inst_core.Inst_controller.n7851\ : std_logic;
signal \Inst_core.Inst_controller.n7852\ : std_logic;
signal \Inst_core.Inst_controller.counter_8\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \Inst_core.Inst_controller.counter_9\ : std_logic;
signal \Inst_core.Inst_controller.n7853\ : std_logic;
signal \Inst_core.Inst_controller.counter_10\ : std_logic;
signal \Inst_core.Inst_controller.n7854\ : std_logic;
signal \Inst_core.Inst_controller.counter_11\ : std_logic;
signal \Inst_core.Inst_controller.n7855\ : std_logic;
signal \Inst_core.Inst_controller.counter_12\ : std_logic;
signal \Inst_core.Inst_controller.n7856\ : std_logic;
signal \Inst_core.Inst_controller.counter_13\ : std_logic;
signal \Inst_core.Inst_controller.n7857\ : std_logic;
signal \Inst_core.Inst_controller.counter_14\ : std_logic;
signal \Inst_core.Inst_controller.n7858\ : std_logic;
signal \Inst_core.Inst_controller.counter_15\ : std_logic;
signal \Inst_core.Inst_controller.n7859\ : std_logic;
signal \Inst_core.Inst_controller.n7860\ : std_logic;
signal \Inst_core.Inst_controller.counter_16\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \Inst_core.Inst_controller.n7861\ : std_logic;
signal \Inst_core.Inst_controller.counter_17\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \xtalClock_c\ : std_logic;
signal \Inst_core.Inst_controller.n3907\ : std_logic;
signal \Inst_core.Inst_controller.n4691\ : std_logic;

signal \xtalClock_wire\ : std_logic;
signal debugleds_wire : std_logic_vector(1 downto 0);
signal input_wire : std_logic_vector(7 downto 0);
signal rx_wire : std_logic;
signal ready50_wire : std_logic;
signal testcnt_wire : std_logic_vector(7 downto 0);
signal tx_wire : std_logic;
signal \GENERIC_FIFO_1.fifo_memory0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \GENERIC_FIFO_1.fifo_memory0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \GENERIC_FIFO_1.fifo_memory0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \GENERIC_FIFO_1.fifo_memory0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \GENERIC_FIFO_1.fifo_memory0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \GENERIC_FIFO_1.fifo_memory1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \GENERIC_FIFO_1.fifo_memory1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \GENERIC_FIFO_1.fifo_memory1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \GENERIC_FIFO_1.fifo_memory1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \GENERIC_FIFO_1.fifo_memory1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \xtalClock_wire\ <= xtalClock;
    debugleds <= debugleds_wire;
    input_wire <= input;
    rx_wire <= rx;
    ready50 <= ready50_wire;
    testcnt <= testcnt_wire;
    tx <= tx_wire;
    outputdata_7 <= \GENERIC_FIFO_1.fifo_memory0_physical_RDATA_wire\(13);
    outputdata_6 <= \GENERIC_FIFO_1.fifo_memory0_physical_RDATA_wire\(9);
    outputdata_5 <= \GENERIC_FIFO_1.fifo_memory0_physical_RDATA_wire\(5);
    outputdata_4 <= \GENERIC_FIFO_1.fifo_memory0_physical_RDATA_wire\(1);
    \GENERIC_FIFO_1.fifo_memory0_physical_RADDR_wire\ <= '0'&\N__15362\&\N__15761\&\N__15782\&\N__16367\&\N__16394\&\N__16409\&\N__16424\&\N__16439\&\N__15887\&\N__15257\;
    \GENERIC_FIFO_1.fifo_memory0_physical_WADDR_wire\ <= '0'&\N__14627\&\N__14672\&\N__14579\&\N__17120\&\N__14879\&\N__14948\&\N__16487\&\N__16535\&\N__16583\&\N__16634\;
    \GENERIC_FIFO_1.fifo_memory0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \GENERIC_FIFO_1.fifo_memory0_physical_WDATA_wire\ <= '0'&'0'&\N__23046\&'0'&'0'&'0'&\N__30462\&'0'&'0'&'0'&\N__25513\&'0'&'0'&'0'&\N__28076\&'0';
    outputdata_3 <= \GENERIC_FIFO_1.fifo_memory1_physical_RDATA_wire\(13);
    outputdata_2 <= \GENERIC_FIFO_1.fifo_memory1_physical_RDATA_wire\(9);
    outputdata_1 <= \GENERIC_FIFO_1.fifo_memory1_physical_RDATA_wire\(5);
    outputdata_0 <= \GENERIC_FIFO_1.fifo_memory1_physical_RDATA_wire\(1);
    \GENERIC_FIFO_1.fifo_memory1_physical_RADDR_wire\ <= '0'&\N__15356\&\N__15755\&\N__15776\&\N__16361\&\N__16388\&\N__16403\&\N__16418\&\N__16433\&\N__15881\&\N__15251\;
    \GENERIC_FIFO_1.fifo_memory1_physical_WADDR_wire\ <= '0'&\N__14621\&\N__14666\&\N__14573\&\N__17112\&\N__14872\&\N__14942\&\N__16479\&\N__16527\&\N__16576\&\N__16626\;
    \GENERIC_FIFO_1.fifo_memory1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \GENERIC_FIFO_1.fifo_memory1_physical_WDATA_wire\ <= '0'&'0'&\N__32337\&'0'&'0'&'0'&\N__30935\&'0'&'0'&'0'&\N__33651\&'0'&'0'&'0'&\N__31817\&'0';

    \GENERIC_FIFO_1.fifo_memory0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \GENERIC_FIFO_1.fifo_memory0_physical_RDATA_wire\,
            RADDR => \GENERIC_FIFO_1.fifo_memory0_physical_RADDR_wire\,
            WADDR => \GENERIC_FIFO_1.fifo_memory0_physical_WADDR_wire\,
            MASK => \GENERIC_FIFO_1.fifo_memory0_physical_MASK_wire\,
            WDATA => \GENERIC_FIFO_1.fifo_memory0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__37486\,
            RE => \N__17350\,
            WCLKE => 'H',
            WCLK => \N__37487\,
            WE => \N__14992\
        );

    \GENERIC_FIFO_1.fifo_memory1_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \GENERIC_FIFO_1.fifo_memory1_physical_RDATA_wire\,
            RADDR => \GENERIC_FIFO_1.fifo_memory1_physical_RADDR_wire\,
            WADDR => \GENERIC_FIFO_1.fifo_memory1_physical_WADDR_wire\,
            MASK => \GENERIC_FIFO_1.fifo_memory1_physical_MASK_wire\,
            WDATA => \GENERIC_FIFO_1.fifo_memory1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__37500\,
            RE => \N__17354\,
            WCLKE => 'H',
            WCLK => \N__37499\,
            WE => \N__14991\
        );

    \xtalClock_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__38004\,
            GLOBALBUFFEROUTPUT => \xtalClock_c\
        );

    \xtalClock_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38006\,
            DIN => \N__38005\,
            DOUT => \N__38004\,
            PACKAGEPIN => \xtalClock_wire\
        );

    \xtalClock_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38006\,
            PADOUT => \N__38005\,
            PADIN => \N__38004\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debugleds_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37995\,
            DIN => \N__37994\,
            DOUT => \N__37993\,
            PACKAGEPIN => debugleds_wire(0)
        );

    \debugleds_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37995\,
            PADOUT => \N__37994\,
            PADIN => \N__37993\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36737\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debugleds_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37986\,
            DIN => \N__37985\,
            DOUT => \N__37984\,
            PACKAGEPIN => debugleds_wire(1)
        );

    \debugleds_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37986\,
            PADOUT => \N__37985\,
            PADIN => \N__37984\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30155\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37977\,
            DIN => \N__37976\,
            DOUT => \N__37975\,
            PACKAGEPIN => input_wire(0)
        );

    \input_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37977\,
            PADOUT => \N__37976\,
            PADIN => \N__37975\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37968\,
            DIN => \N__37967\,
            DOUT => \N__37966\,
            PACKAGEPIN => input_wire(1)
        );

    \input_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37968\,
            PADOUT => \N__37967\,
            PADIN => \N__37966\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37959\,
            DIN => \N__37958\,
            DOUT => \N__37957\,
            PACKAGEPIN => input_wire(2)
        );

    \input_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37959\,
            PADOUT => \N__37958\,
            PADIN => \N__37957\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37950\,
            DIN => \N__37949\,
            DOUT => \N__37948\,
            PACKAGEPIN => input_wire(3)
        );

    \input_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37950\,
            PADOUT => \N__37949\,
            PADIN => \N__37948\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37941\,
            DIN => \N__37940\,
            DOUT => \N__37939\,
            PACKAGEPIN => input_wire(4)
        );

    \input_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37941\,
            PADOUT => \N__37940\,
            PADIN => \N__37939\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37932\,
            DIN => \N__37931\,
            DOUT => \N__37930\,
            PACKAGEPIN => input_wire(5)
        );

    \input_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37932\,
            PADOUT => \N__37931\,
            PADIN => \N__37930\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37923\,
            DIN => \N__37922\,
            DOUT => \N__37921\,
            PACKAGEPIN => input_wire(6)
        );

    \input_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37923\,
            PADOUT => \N__37922\,
            PADIN => \N__37921\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \input_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37914\,
            DIN => \N__37913\,
            DOUT => \N__37912\,
            PACKAGEPIN => input_wire(7)
        );

    \input_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37914\,
            PADOUT => \N__37913\,
            PADIN => \N__37912\,
            CLOCKENABLE => 'H',
            DIN0 => input_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \nstate_2__N_139_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37905\,
            DIN => \N__37904\,
            DOUT => \N__37903\,
            PACKAGEPIN => rx_wire
        );

    \nstate_2__N_139_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37905\,
            PADOUT => \N__37904\,
            PADIN => \N__37903\,
            CLOCKENABLE => 'H',
            DIN0 => \nstate_2__N_139_c_1\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ready50_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37896\,
            DIN => \N__37895\,
            DOUT => \N__37894\,
            PACKAGEPIN => ready50_wire
        );

    \ready50_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37896\,
            PADOUT => \N__37895\,
            PADIN => \N__37894\,
            CLOCKENABLE => \N__32228\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31956\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__37621\,
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37887\,
            DIN => \N__37886\,
            DOUT => \N__37885\,
            PACKAGEPIN => testcnt_wire(0)
        );

    \testcnt_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37887\,
            PADOUT => \N__37886\,
            PADIN => \N__37885\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19487\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37878\,
            DIN => \N__37877\,
            DOUT => \N__37876\,
            PACKAGEPIN => testcnt_wire(1)
        );

    \testcnt_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37878\,
            PADOUT => \N__37877\,
            PADIN => \N__37876\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19910\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37869\,
            DIN => \N__37868\,
            DOUT => \N__37867\,
            PACKAGEPIN => testcnt_wire(2)
        );

    \testcnt_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37869\,
            PADOUT => \N__37868\,
            PADIN => \N__37867\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19889\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37860\,
            DIN => \N__37859\,
            DOUT => \N__37858\,
            PACKAGEPIN => testcnt_wire(3)
        );

    \testcnt_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37860\,
            PADOUT => \N__37859\,
            PADIN => \N__37858\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19868\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37851\,
            DIN => \N__37850\,
            DOUT => \N__37849\,
            PACKAGEPIN => testcnt_wire(4)
        );

    \testcnt_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37851\,
            PADOUT => \N__37850\,
            PADIN => \N__37849\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19853\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37842\,
            DIN => \N__37841\,
            DOUT => \N__37840\,
            PACKAGEPIN => testcnt_wire(5)
        );

    \testcnt_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37842\,
            PADOUT => \N__37841\,
            PADIN => \N__37840\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19838\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37833\,
            DIN => \N__37832\,
            DOUT => \N__37831\,
            PACKAGEPIN => testcnt_wire(6)
        );

    \testcnt_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37833\,
            PADOUT => \N__37832\,
            PADIN => \N__37831\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19823\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \testcnt_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37824\,
            DIN => \N__37823\,
            DOUT => \N__37822\,
            PACKAGEPIN => testcnt_wire(7)
        );

    \testcnt_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37824\,
            PADOUT => \N__37823\,
            PADIN => \N__37822\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19799\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37815\,
            DIN => \N__37814\,
            DOUT => \N__37813\,
            PACKAGEPIN => tx_wire
        );

    \tx_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37815\,
            PADOUT => \N__37814\,
            PADIN => \N__37813\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13559\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__9296\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37790\
        );

    \I__9295\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37790\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__37790\,
            I => \N__37786\
        );

    \I__9293\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37783\
        );

    \I__9292\ : Span4Mux_h
    port map (
            O => \N__37786\,
            I => \N__37780\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__37783\,
            I => \Inst_core.Inst_controller.counter_12\
        );

    \I__9290\ : Odrv4
    port map (
            O => \N__37780\,
            I => \Inst_core.Inst_controller.counter_12\
        );

    \I__9289\ : InMux
    port map (
            O => \N__37775\,
            I => \Inst_core.Inst_controller.n7856\
        );

    \I__9288\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37766\
        );

    \I__9287\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37766\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__37766\,
            I => \N__37762\
        );

    \I__9285\ : InMux
    port map (
            O => \N__37765\,
            I => \N__37759\
        );

    \I__9284\ : Span4Mux_v
    port map (
            O => \N__37762\,
            I => \N__37756\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__37759\,
            I => \Inst_core.Inst_controller.counter_13\
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__37756\,
            I => \Inst_core.Inst_controller.counter_13\
        );

    \I__9281\ : InMux
    port map (
            O => \N__37751\,
            I => \Inst_core.Inst_controller.n7857\
        );

    \I__9280\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37742\
        );

    \I__9279\ : InMux
    port map (
            O => \N__37747\,
            I => \N__37742\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__37742\,
            I => \N__37738\
        );

    \I__9277\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37735\
        );

    \I__9276\ : Span4Mux_h
    port map (
            O => \N__37738\,
            I => \N__37732\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__37735\,
            I => \Inst_core.Inst_controller.counter_14\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__37732\,
            I => \Inst_core.Inst_controller.counter_14\
        );

    \I__9273\ : InMux
    port map (
            O => \N__37727\,
            I => \Inst_core.Inst_controller.n7858\
        );

    \I__9272\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37720\
        );

    \I__9271\ : InMux
    port map (
            O => \N__37723\,
            I => \N__37716\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__37720\,
            I => \N__37713\
        );

    \I__9269\ : InMux
    port map (
            O => \N__37719\,
            I => \N__37710\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37705\
        );

    \I__9267\ : Span4Mux_h
    port map (
            O => \N__37713\,
            I => \N__37705\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__37710\,
            I => \Inst_core.Inst_controller.counter_15\
        );

    \I__9265\ : Odrv4
    port map (
            O => \N__37705\,
            I => \Inst_core.Inst_controller.counter_15\
        );

    \I__9264\ : InMux
    port map (
            O => \N__37700\,
            I => \Inst_core.Inst_controller.n7859\
        );

    \I__9263\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37693\
        );

    \I__9262\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37690\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__37693\,
            I => \N__37687\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__37690\,
            I => \N__37681\
        );

    \I__9259\ : Span4Mux_h
    port map (
            O => \N__37687\,
            I => \N__37681\
        );

    \I__9258\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37678\
        );

    \I__9257\ : Span4Mux_h
    port map (
            O => \N__37681\,
            I => \N__37675\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__37678\,
            I => \Inst_core.Inst_controller.counter_16\
        );

    \I__9255\ : Odrv4
    port map (
            O => \N__37675\,
            I => \Inst_core.Inst_controller.counter_16\
        );

    \I__9254\ : InMux
    port map (
            O => \N__37670\,
            I => \bfn_12_14_0_\
        );

    \I__9253\ : InMux
    port map (
            O => \N__37667\,
            I => \Inst_core.Inst_controller.n7861\
        );

    \I__9252\ : InMux
    port map (
            O => \N__37664\,
            I => \N__37660\
        );

    \I__9251\ : InMux
    port map (
            O => \N__37663\,
            I => \N__37657\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__37660\,
            I => \N__37653\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__37657\,
            I => \N__37650\
        );

    \I__9248\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37647\
        );

    \I__9247\ : Span4Mux_h
    port map (
            O => \N__37653\,
            I => \N__37644\
        );

    \I__9246\ : Span4Mux_h
    port map (
            O => \N__37650\,
            I => \N__37641\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__37647\,
            I => \N__37636\
        );

    \I__9244\ : Span4Mux_v
    port map (
            O => \N__37644\,
            I => \N__37636\
        );

    \I__9243\ : Span4Mux_h
    port map (
            O => \N__37641\,
            I => \N__37633\
        );

    \I__9242\ : Odrv4
    port map (
            O => \N__37636\,
            I => \Inst_core.Inst_controller.counter_17\
        );

    \I__9241\ : Odrv4
    port map (
            O => \N__37633\,
            I => \Inst_core.Inst_controller.counter_17\
        );

    \I__9240\ : ClkMux
    port map (
            O => \N__37628\,
            I => \N__37163\
        );

    \I__9239\ : ClkMux
    port map (
            O => \N__37627\,
            I => \N__37163\
        );

    \I__9238\ : ClkMux
    port map (
            O => \N__37626\,
            I => \N__37163\
        );

    \I__9237\ : ClkMux
    port map (
            O => \N__37625\,
            I => \N__37163\
        );

    \I__9236\ : ClkMux
    port map (
            O => \N__37624\,
            I => \N__37163\
        );

    \I__9235\ : ClkMux
    port map (
            O => \N__37623\,
            I => \N__37163\
        );

    \I__9234\ : ClkMux
    port map (
            O => \N__37622\,
            I => \N__37163\
        );

    \I__9233\ : ClkMux
    port map (
            O => \N__37621\,
            I => \N__37163\
        );

    \I__9232\ : ClkMux
    port map (
            O => \N__37620\,
            I => \N__37163\
        );

    \I__9231\ : ClkMux
    port map (
            O => \N__37619\,
            I => \N__37163\
        );

    \I__9230\ : ClkMux
    port map (
            O => \N__37618\,
            I => \N__37163\
        );

    \I__9229\ : ClkMux
    port map (
            O => \N__37617\,
            I => \N__37163\
        );

    \I__9228\ : ClkMux
    port map (
            O => \N__37616\,
            I => \N__37163\
        );

    \I__9227\ : ClkMux
    port map (
            O => \N__37615\,
            I => \N__37163\
        );

    \I__9226\ : ClkMux
    port map (
            O => \N__37614\,
            I => \N__37163\
        );

    \I__9225\ : ClkMux
    port map (
            O => \N__37613\,
            I => \N__37163\
        );

    \I__9224\ : ClkMux
    port map (
            O => \N__37612\,
            I => \N__37163\
        );

    \I__9223\ : ClkMux
    port map (
            O => \N__37611\,
            I => \N__37163\
        );

    \I__9222\ : ClkMux
    port map (
            O => \N__37610\,
            I => \N__37163\
        );

    \I__9221\ : ClkMux
    port map (
            O => \N__37609\,
            I => \N__37163\
        );

    \I__9220\ : ClkMux
    port map (
            O => \N__37608\,
            I => \N__37163\
        );

    \I__9219\ : ClkMux
    port map (
            O => \N__37607\,
            I => \N__37163\
        );

    \I__9218\ : ClkMux
    port map (
            O => \N__37606\,
            I => \N__37163\
        );

    \I__9217\ : ClkMux
    port map (
            O => \N__37605\,
            I => \N__37163\
        );

    \I__9216\ : ClkMux
    port map (
            O => \N__37604\,
            I => \N__37163\
        );

    \I__9215\ : ClkMux
    port map (
            O => \N__37603\,
            I => \N__37163\
        );

    \I__9214\ : ClkMux
    port map (
            O => \N__37602\,
            I => \N__37163\
        );

    \I__9213\ : ClkMux
    port map (
            O => \N__37601\,
            I => \N__37163\
        );

    \I__9212\ : ClkMux
    port map (
            O => \N__37600\,
            I => \N__37163\
        );

    \I__9211\ : ClkMux
    port map (
            O => \N__37599\,
            I => \N__37163\
        );

    \I__9210\ : ClkMux
    port map (
            O => \N__37598\,
            I => \N__37163\
        );

    \I__9209\ : ClkMux
    port map (
            O => \N__37597\,
            I => \N__37163\
        );

    \I__9208\ : ClkMux
    port map (
            O => \N__37596\,
            I => \N__37163\
        );

    \I__9207\ : ClkMux
    port map (
            O => \N__37595\,
            I => \N__37163\
        );

    \I__9206\ : ClkMux
    port map (
            O => \N__37594\,
            I => \N__37163\
        );

    \I__9205\ : ClkMux
    port map (
            O => \N__37593\,
            I => \N__37163\
        );

    \I__9204\ : ClkMux
    port map (
            O => \N__37592\,
            I => \N__37163\
        );

    \I__9203\ : ClkMux
    port map (
            O => \N__37591\,
            I => \N__37163\
        );

    \I__9202\ : ClkMux
    port map (
            O => \N__37590\,
            I => \N__37163\
        );

    \I__9201\ : ClkMux
    port map (
            O => \N__37589\,
            I => \N__37163\
        );

    \I__9200\ : ClkMux
    port map (
            O => \N__37588\,
            I => \N__37163\
        );

    \I__9199\ : ClkMux
    port map (
            O => \N__37587\,
            I => \N__37163\
        );

    \I__9198\ : ClkMux
    port map (
            O => \N__37586\,
            I => \N__37163\
        );

    \I__9197\ : ClkMux
    port map (
            O => \N__37585\,
            I => \N__37163\
        );

    \I__9196\ : ClkMux
    port map (
            O => \N__37584\,
            I => \N__37163\
        );

    \I__9195\ : ClkMux
    port map (
            O => \N__37583\,
            I => \N__37163\
        );

    \I__9194\ : ClkMux
    port map (
            O => \N__37582\,
            I => \N__37163\
        );

    \I__9193\ : ClkMux
    port map (
            O => \N__37581\,
            I => \N__37163\
        );

    \I__9192\ : ClkMux
    port map (
            O => \N__37580\,
            I => \N__37163\
        );

    \I__9191\ : ClkMux
    port map (
            O => \N__37579\,
            I => \N__37163\
        );

    \I__9190\ : ClkMux
    port map (
            O => \N__37578\,
            I => \N__37163\
        );

    \I__9189\ : ClkMux
    port map (
            O => \N__37577\,
            I => \N__37163\
        );

    \I__9188\ : ClkMux
    port map (
            O => \N__37576\,
            I => \N__37163\
        );

    \I__9187\ : ClkMux
    port map (
            O => \N__37575\,
            I => \N__37163\
        );

    \I__9186\ : ClkMux
    port map (
            O => \N__37574\,
            I => \N__37163\
        );

    \I__9185\ : ClkMux
    port map (
            O => \N__37573\,
            I => \N__37163\
        );

    \I__9184\ : ClkMux
    port map (
            O => \N__37572\,
            I => \N__37163\
        );

    \I__9183\ : ClkMux
    port map (
            O => \N__37571\,
            I => \N__37163\
        );

    \I__9182\ : ClkMux
    port map (
            O => \N__37570\,
            I => \N__37163\
        );

    \I__9181\ : ClkMux
    port map (
            O => \N__37569\,
            I => \N__37163\
        );

    \I__9180\ : ClkMux
    port map (
            O => \N__37568\,
            I => \N__37163\
        );

    \I__9179\ : ClkMux
    port map (
            O => \N__37567\,
            I => \N__37163\
        );

    \I__9178\ : ClkMux
    port map (
            O => \N__37566\,
            I => \N__37163\
        );

    \I__9177\ : ClkMux
    port map (
            O => \N__37565\,
            I => \N__37163\
        );

    \I__9176\ : ClkMux
    port map (
            O => \N__37564\,
            I => \N__37163\
        );

    \I__9175\ : ClkMux
    port map (
            O => \N__37563\,
            I => \N__37163\
        );

    \I__9174\ : ClkMux
    port map (
            O => \N__37562\,
            I => \N__37163\
        );

    \I__9173\ : ClkMux
    port map (
            O => \N__37561\,
            I => \N__37163\
        );

    \I__9172\ : ClkMux
    port map (
            O => \N__37560\,
            I => \N__37163\
        );

    \I__9171\ : ClkMux
    port map (
            O => \N__37559\,
            I => \N__37163\
        );

    \I__9170\ : ClkMux
    port map (
            O => \N__37558\,
            I => \N__37163\
        );

    \I__9169\ : ClkMux
    port map (
            O => \N__37557\,
            I => \N__37163\
        );

    \I__9168\ : ClkMux
    port map (
            O => \N__37556\,
            I => \N__37163\
        );

    \I__9167\ : ClkMux
    port map (
            O => \N__37555\,
            I => \N__37163\
        );

    \I__9166\ : ClkMux
    port map (
            O => \N__37554\,
            I => \N__37163\
        );

    \I__9165\ : ClkMux
    port map (
            O => \N__37553\,
            I => \N__37163\
        );

    \I__9164\ : ClkMux
    port map (
            O => \N__37552\,
            I => \N__37163\
        );

    \I__9163\ : ClkMux
    port map (
            O => \N__37551\,
            I => \N__37163\
        );

    \I__9162\ : ClkMux
    port map (
            O => \N__37550\,
            I => \N__37163\
        );

    \I__9161\ : ClkMux
    port map (
            O => \N__37549\,
            I => \N__37163\
        );

    \I__9160\ : ClkMux
    port map (
            O => \N__37548\,
            I => \N__37163\
        );

    \I__9159\ : ClkMux
    port map (
            O => \N__37547\,
            I => \N__37163\
        );

    \I__9158\ : ClkMux
    port map (
            O => \N__37546\,
            I => \N__37163\
        );

    \I__9157\ : ClkMux
    port map (
            O => \N__37545\,
            I => \N__37163\
        );

    \I__9156\ : ClkMux
    port map (
            O => \N__37544\,
            I => \N__37163\
        );

    \I__9155\ : ClkMux
    port map (
            O => \N__37543\,
            I => \N__37163\
        );

    \I__9154\ : ClkMux
    port map (
            O => \N__37542\,
            I => \N__37163\
        );

    \I__9153\ : ClkMux
    port map (
            O => \N__37541\,
            I => \N__37163\
        );

    \I__9152\ : ClkMux
    port map (
            O => \N__37540\,
            I => \N__37163\
        );

    \I__9151\ : ClkMux
    port map (
            O => \N__37539\,
            I => \N__37163\
        );

    \I__9150\ : ClkMux
    port map (
            O => \N__37538\,
            I => \N__37163\
        );

    \I__9149\ : ClkMux
    port map (
            O => \N__37537\,
            I => \N__37163\
        );

    \I__9148\ : ClkMux
    port map (
            O => \N__37536\,
            I => \N__37163\
        );

    \I__9147\ : ClkMux
    port map (
            O => \N__37535\,
            I => \N__37163\
        );

    \I__9146\ : ClkMux
    port map (
            O => \N__37534\,
            I => \N__37163\
        );

    \I__9145\ : ClkMux
    port map (
            O => \N__37533\,
            I => \N__37163\
        );

    \I__9144\ : ClkMux
    port map (
            O => \N__37532\,
            I => \N__37163\
        );

    \I__9143\ : ClkMux
    port map (
            O => \N__37531\,
            I => \N__37163\
        );

    \I__9142\ : ClkMux
    port map (
            O => \N__37530\,
            I => \N__37163\
        );

    \I__9141\ : ClkMux
    port map (
            O => \N__37529\,
            I => \N__37163\
        );

    \I__9140\ : ClkMux
    port map (
            O => \N__37528\,
            I => \N__37163\
        );

    \I__9139\ : ClkMux
    port map (
            O => \N__37527\,
            I => \N__37163\
        );

    \I__9138\ : ClkMux
    port map (
            O => \N__37526\,
            I => \N__37163\
        );

    \I__9137\ : ClkMux
    port map (
            O => \N__37525\,
            I => \N__37163\
        );

    \I__9136\ : ClkMux
    port map (
            O => \N__37524\,
            I => \N__37163\
        );

    \I__9135\ : ClkMux
    port map (
            O => \N__37523\,
            I => \N__37163\
        );

    \I__9134\ : ClkMux
    port map (
            O => \N__37522\,
            I => \N__37163\
        );

    \I__9133\ : ClkMux
    port map (
            O => \N__37521\,
            I => \N__37163\
        );

    \I__9132\ : ClkMux
    port map (
            O => \N__37520\,
            I => \N__37163\
        );

    \I__9131\ : ClkMux
    port map (
            O => \N__37519\,
            I => \N__37163\
        );

    \I__9130\ : ClkMux
    port map (
            O => \N__37518\,
            I => \N__37163\
        );

    \I__9129\ : ClkMux
    port map (
            O => \N__37517\,
            I => \N__37163\
        );

    \I__9128\ : ClkMux
    port map (
            O => \N__37516\,
            I => \N__37163\
        );

    \I__9127\ : ClkMux
    port map (
            O => \N__37515\,
            I => \N__37163\
        );

    \I__9126\ : ClkMux
    port map (
            O => \N__37514\,
            I => \N__37163\
        );

    \I__9125\ : ClkMux
    port map (
            O => \N__37513\,
            I => \N__37163\
        );

    \I__9124\ : ClkMux
    port map (
            O => \N__37512\,
            I => \N__37163\
        );

    \I__9123\ : ClkMux
    port map (
            O => \N__37511\,
            I => \N__37163\
        );

    \I__9122\ : ClkMux
    port map (
            O => \N__37510\,
            I => \N__37163\
        );

    \I__9121\ : ClkMux
    port map (
            O => \N__37509\,
            I => \N__37163\
        );

    \I__9120\ : ClkMux
    port map (
            O => \N__37508\,
            I => \N__37163\
        );

    \I__9119\ : ClkMux
    port map (
            O => \N__37507\,
            I => \N__37163\
        );

    \I__9118\ : ClkMux
    port map (
            O => \N__37506\,
            I => \N__37163\
        );

    \I__9117\ : ClkMux
    port map (
            O => \N__37505\,
            I => \N__37163\
        );

    \I__9116\ : ClkMux
    port map (
            O => \N__37504\,
            I => \N__37163\
        );

    \I__9115\ : ClkMux
    port map (
            O => \N__37503\,
            I => \N__37163\
        );

    \I__9114\ : ClkMux
    port map (
            O => \N__37502\,
            I => \N__37163\
        );

    \I__9113\ : ClkMux
    port map (
            O => \N__37501\,
            I => \N__37163\
        );

    \I__9112\ : ClkMux
    port map (
            O => \N__37500\,
            I => \N__37163\
        );

    \I__9111\ : ClkMux
    port map (
            O => \N__37499\,
            I => \N__37163\
        );

    \I__9110\ : ClkMux
    port map (
            O => \N__37498\,
            I => \N__37163\
        );

    \I__9109\ : ClkMux
    port map (
            O => \N__37497\,
            I => \N__37163\
        );

    \I__9108\ : ClkMux
    port map (
            O => \N__37496\,
            I => \N__37163\
        );

    \I__9107\ : ClkMux
    port map (
            O => \N__37495\,
            I => \N__37163\
        );

    \I__9106\ : ClkMux
    port map (
            O => \N__37494\,
            I => \N__37163\
        );

    \I__9105\ : ClkMux
    port map (
            O => \N__37493\,
            I => \N__37163\
        );

    \I__9104\ : ClkMux
    port map (
            O => \N__37492\,
            I => \N__37163\
        );

    \I__9103\ : ClkMux
    port map (
            O => \N__37491\,
            I => \N__37163\
        );

    \I__9102\ : ClkMux
    port map (
            O => \N__37490\,
            I => \N__37163\
        );

    \I__9101\ : ClkMux
    port map (
            O => \N__37489\,
            I => \N__37163\
        );

    \I__9100\ : ClkMux
    port map (
            O => \N__37488\,
            I => \N__37163\
        );

    \I__9099\ : ClkMux
    port map (
            O => \N__37487\,
            I => \N__37163\
        );

    \I__9098\ : ClkMux
    port map (
            O => \N__37486\,
            I => \N__37163\
        );

    \I__9097\ : ClkMux
    port map (
            O => \N__37485\,
            I => \N__37163\
        );

    \I__9096\ : ClkMux
    port map (
            O => \N__37484\,
            I => \N__37163\
        );

    \I__9095\ : ClkMux
    port map (
            O => \N__37483\,
            I => \N__37163\
        );

    \I__9094\ : ClkMux
    port map (
            O => \N__37482\,
            I => \N__37163\
        );

    \I__9093\ : ClkMux
    port map (
            O => \N__37481\,
            I => \N__37163\
        );

    \I__9092\ : ClkMux
    port map (
            O => \N__37480\,
            I => \N__37163\
        );

    \I__9091\ : ClkMux
    port map (
            O => \N__37479\,
            I => \N__37163\
        );

    \I__9090\ : ClkMux
    port map (
            O => \N__37478\,
            I => \N__37163\
        );

    \I__9089\ : ClkMux
    port map (
            O => \N__37477\,
            I => \N__37163\
        );

    \I__9088\ : ClkMux
    port map (
            O => \N__37476\,
            I => \N__37163\
        );

    \I__9087\ : ClkMux
    port map (
            O => \N__37475\,
            I => \N__37163\
        );

    \I__9086\ : ClkMux
    port map (
            O => \N__37474\,
            I => \N__37163\
        );

    \I__9085\ : GlobalMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__9084\ : gio2CtrlBuf
    port map (
            O => \N__37160\,
            I => \xtalClock_c\
        );

    \I__9083\ : CEMux
    port map (
            O => \N__37157\,
            I => \N__37153\
        );

    \I__9082\ : CEMux
    port map (
            O => \N__37156\,
            I => \N__37149\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__37153\,
            I => \N__37146\
        );

    \I__9080\ : CEMux
    port map (
            O => \N__37152\,
            I => \N__37143\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__37149\,
            I => \N__37140\
        );

    \I__9078\ : Span4Mux_s0_h
    port map (
            O => \N__37146\,
            I => \N__37135\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__37143\,
            I => \N__37135\
        );

    \I__9076\ : Span4Mux_v
    port map (
            O => \N__37140\,
            I => \N__37132\
        );

    \I__9075\ : Span4Mux_v
    port map (
            O => \N__37135\,
            I => \N__37127\
        );

    \I__9074\ : Span4Mux_s0_h
    port map (
            O => \N__37132\,
            I => \N__37127\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__37127\,
            I => \Inst_core.Inst_controller.n3907\
        );

    \I__9072\ : SRMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__9070\ : Span4Mux_s1_h
    port map (
            O => \N__37118\,
            I => \N__37113\
        );

    \I__9069\ : SRMux
    port map (
            O => \N__37117\,
            I => \N__37110\
        );

    \I__9068\ : SRMux
    port map (
            O => \N__37116\,
            I => \N__37107\
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__37113\,
            I => \Inst_core.Inst_controller.n4691\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__37110\,
            I => \Inst_core.Inst_controller.n4691\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__37107\,
            I => \Inst_core.Inst_controller.n4691\
        );

    \I__9064\ : InMux
    port map (
            O => \N__37100\,
            I => \N__37095\
        );

    \I__9063\ : InMux
    port map (
            O => \N__37099\,
            I => \N__37092\
        );

    \I__9062\ : InMux
    port map (
            O => \N__37098\,
            I => \N__37089\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__37095\,
            I => \Inst_core.Inst_controller.counter_4\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__37092\,
            I => \Inst_core.Inst_controller.counter_4\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__37089\,
            I => \Inst_core.Inst_controller.counter_4\
        );

    \I__9058\ : InMux
    port map (
            O => \N__37082\,
            I => \Inst_core.Inst_controller.n7848\
        );

    \I__9057\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37075\
        );

    \I__9056\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37072\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__37075\,
            I => \N__37066\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__37072\,
            I => \N__37066\
        );

    \I__9053\ : InMux
    port map (
            O => \N__37071\,
            I => \N__37063\
        );

    \I__9052\ : Span4Mux_h
    port map (
            O => \N__37066\,
            I => \N__37060\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__37063\,
            I => \Inst_core.Inst_controller.counter_5\
        );

    \I__9050\ : Odrv4
    port map (
            O => \N__37060\,
            I => \Inst_core.Inst_controller.counter_5\
        );

    \I__9049\ : InMux
    port map (
            O => \N__37055\,
            I => \Inst_core.Inst_controller.n7849\
        );

    \I__9048\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37048\
        );

    \I__9047\ : InMux
    port map (
            O => \N__37051\,
            I => \N__37045\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__37048\,
            I => \N__37039\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__37045\,
            I => \N__37039\
        );

    \I__9044\ : InMux
    port map (
            O => \N__37044\,
            I => \N__37036\
        );

    \I__9043\ : Span4Mux_h
    port map (
            O => \N__37039\,
            I => \N__37033\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__37036\,
            I => \Inst_core.Inst_controller.counter_6\
        );

    \I__9041\ : Odrv4
    port map (
            O => \N__37033\,
            I => \Inst_core.Inst_controller.counter_6\
        );

    \I__9040\ : InMux
    port map (
            O => \N__37028\,
            I => \Inst_core.Inst_controller.n7850\
        );

    \I__9039\ : InMux
    port map (
            O => \N__37025\,
            I => \N__37021\
        );

    \I__9038\ : InMux
    port map (
            O => \N__37024\,
            I => \N__37018\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__37021\,
            I => \N__37015\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__37018\,
            I => \N__37011\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__37015\,
            I => \N__37008\
        );

    \I__9034\ : InMux
    port map (
            O => \N__37014\,
            I => \N__37005\
        );

    \I__9033\ : Span4Mux_v
    port map (
            O => \N__37011\,
            I => \N__37002\
        );

    \I__9032\ : Span4Mux_h
    port map (
            O => \N__37008\,
            I => \N__36999\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__37005\,
            I => \Inst_core.Inst_controller.counter_7\
        );

    \I__9030\ : Odrv4
    port map (
            O => \N__37002\,
            I => \Inst_core.Inst_controller.counter_7\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__36999\,
            I => \Inst_core.Inst_controller.counter_7\
        );

    \I__9028\ : InMux
    port map (
            O => \N__36992\,
            I => \Inst_core.Inst_controller.n7851\
        );

    \I__9027\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36985\
        );

    \I__9026\ : InMux
    port map (
            O => \N__36988\,
            I => \N__36982\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__36985\,
            I => \N__36979\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__36982\,
            I => \N__36975\
        );

    \I__9023\ : Span4Mux_h
    port map (
            O => \N__36979\,
            I => \N__36972\
        );

    \I__9022\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36969\
        );

    \I__9021\ : Span4Mux_h
    port map (
            O => \N__36975\,
            I => \N__36966\
        );

    \I__9020\ : Span4Mux_h
    port map (
            O => \N__36972\,
            I => \N__36963\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__36969\,
            I => \Inst_core.Inst_controller.counter_8\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__36966\,
            I => \Inst_core.Inst_controller.counter_8\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__36963\,
            I => \Inst_core.Inst_controller.counter_8\
        );

    \I__9016\ : InMux
    port map (
            O => \N__36956\,
            I => \bfn_12_13_0_\
        );

    \I__9015\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36947\
        );

    \I__9014\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36947\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__36947\,
            I => \N__36943\
        );

    \I__9012\ : InMux
    port map (
            O => \N__36946\,
            I => \N__36940\
        );

    \I__9011\ : Span4Mux_h
    port map (
            O => \N__36943\,
            I => \N__36937\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__36940\,
            I => \Inst_core.Inst_controller.counter_9\
        );

    \I__9009\ : Odrv4
    port map (
            O => \N__36937\,
            I => \Inst_core.Inst_controller.counter_9\
        );

    \I__9008\ : InMux
    port map (
            O => \N__36932\,
            I => \Inst_core.Inst_controller.n7853\
        );

    \I__9007\ : InMux
    port map (
            O => \N__36929\,
            I => \N__36925\
        );

    \I__9006\ : InMux
    port map (
            O => \N__36928\,
            I => \N__36922\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__36925\,
            I => \N__36916\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__36922\,
            I => \N__36916\
        );

    \I__9003\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36913\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__36916\,
            I => \N__36910\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__36913\,
            I => \Inst_core.Inst_controller.counter_10\
        );

    \I__9000\ : Odrv4
    port map (
            O => \N__36910\,
            I => \Inst_core.Inst_controller.counter_10\
        );

    \I__8999\ : InMux
    port map (
            O => \N__36905\,
            I => \Inst_core.Inst_controller.n7854\
        );

    \I__8998\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36898\
        );

    \I__8997\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36895\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__36898\,
            I => \N__36889\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__36895\,
            I => \N__36889\
        );

    \I__8994\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36886\
        );

    \I__8993\ : Span4Mux_h
    port map (
            O => \N__36889\,
            I => \N__36883\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__36886\,
            I => \Inst_core.Inst_controller.counter_11\
        );

    \I__8991\ : Odrv4
    port map (
            O => \N__36883\,
            I => \Inst_core.Inst_controller.counter_11\
        );

    \I__8990\ : InMux
    port map (
            O => \N__36878\,
            I => \Inst_core.Inst_controller.n7855\
        );

    \I__8989\ : SRMux
    port map (
            O => \N__36875\,
            I => \N__36868\
        );

    \I__8988\ : CascadeMux
    port map (
            O => \N__36874\,
            I => \N__36861\
        );

    \I__8987\ : CascadeMux
    port map (
            O => \N__36873\,
            I => \N__36855\
        );

    \I__8986\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36851\
        );

    \I__8985\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36848\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36845\
        );

    \I__8983\ : CascadeMux
    port map (
            O => \N__36867\,
            I => \N__36841\
        );

    \I__8982\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36838\
        );

    \I__8981\ : SRMux
    port map (
            O => \N__36865\,
            I => \N__36835\
        );

    \I__8980\ : SRMux
    port map (
            O => \N__36864\,
            I => \N__36832\
        );

    \I__8979\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36823\
        );

    \I__8978\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36823\
        );

    \I__8977\ : InMux
    port map (
            O => \N__36859\,
            I => \N__36823\
        );

    \I__8976\ : InMux
    port map (
            O => \N__36858\,
            I => \N__36823\
        );

    \I__8975\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36818\
        );

    \I__8974\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36818\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__36851\,
            I => \N__36813\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__36848\,
            I => \N__36813\
        );

    \I__8971\ : Span4Mux_v
    port map (
            O => \N__36845\,
            I => \N__36809\
        );

    \I__8970\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36803\
        );

    \I__8969\ : InMux
    port map (
            O => \N__36841\,
            I => \N__36803\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__36838\,
            I => \N__36800\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__36835\,
            I => \N__36797\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__36832\,
            I => \N__36790\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__36823\,
            I => \N__36790\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__36818\,
            I => \N__36790\
        );

    \I__8963\ : Span4Mux_s3_h
    port map (
            O => \N__36813\,
            I => \N__36787\
        );

    \I__8962\ : InMux
    port map (
            O => \N__36812\,
            I => \N__36784\
        );

    \I__8961\ : Span4Mux_h
    port map (
            O => \N__36809\,
            I => \N__36781\
        );

    \I__8960\ : InMux
    port map (
            O => \N__36808\,
            I => \N__36778\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__36803\,
            I => \N__36773\
        );

    \I__8958\ : Sp12to4
    port map (
            O => \N__36800\,
            I => \N__36773\
        );

    \I__8957\ : Span4Mux_s3_v
    port map (
            O => \N__36797\,
            I => \N__36770\
        );

    \I__8956\ : Span4Mux_s3_v
    port map (
            O => \N__36790\,
            I => \N__36767\
        );

    \I__8955\ : Span4Mux_h
    port map (
            O => \N__36787\,
            I => \N__36762\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__36784\,
            I => \N__36762\
        );

    \I__8953\ : Span4Mux_h
    port map (
            O => \N__36781\,
            I => \N__36759\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__36778\,
            I => \N__36756\
        );

    \I__8951\ : Span12Mux_s8_h
    port map (
            O => \N__36773\,
            I => \N__36753\
        );

    \I__8950\ : Span4Mux_h
    port map (
            O => \N__36770\,
            I => \N__36746\
        );

    \I__8949\ : Span4Mux_h
    port map (
            O => \N__36767\,
            I => \N__36746\
        );

    \I__8948\ : Span4Mux_v
    port map (
            O => \N__36762\,
            I => \N__36746\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__36759\,
            I => \Inst_core.resetCmd\
        );

    \I__8946\ : Odrv12
    port map (
            O => \N__36756\,
            I => \Inst_core.resetCmd\
        );

    \I__8945\ : Odrv12
    port map (
            O => \N__36753\,
            I => \Inst_core.resetCmd\
        );

    \I__8944\ : Odrv4
    port map (
            O => \N__36746\,
            I => \Inst_core.resetCmd\
        );

    \I__8943\ : IoInMux
    port map (
            O => \N__36737\,
            I => \N__36734\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__36734\,
            I => debugleds_c_0
        );

    \I__8941\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36725\
        );

    \I__8940\ : InMux
    port map (
            O => \N__36730\,
            I => \N__36725\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__8938\ : Span12Mux_s0_h
    port map (
            O => \N__36722\,
            I => \N__36719\
        );

    \I__8937\ : Odrv12
    port map (
            O => \N__36719\,
            I => busy
        );

    \I__8936\ : CascadeMux
    port map (
            O => \N__36716\,
            I => \N__36713\
        );

    \I__8935\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__36710\,
            I => \Inst_core.Inst_controller.nstate_1_N_825_0\
        );

    \I__8933\ : CascadeMux
    port map (
            O => \N__36707\,
            I => \N__36702\
        );

    \I__8932\ : InMux
    port map (
            O => \N__36706\,
            I => \N__36692\
        );

    \I__8931\ : InMux
    port map (
            O => \N__36705\,
            I => \N__36692\
        );

    \I__8930\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36692\
        );

    \I__8929\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36692\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__36692\,
            I => \Inst_core.Inst_controller.n320\
        );

    \I__8927\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36680\
        );

    \I__8926\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36680\
        );

    \I__8925\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36680\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__36680\,
            I => \N__36677\
        );

    \I__8923\ : Odrv12
    port map (
            O => \N__36677\,
            I => \Inst_core.Inst_controller.nstate_1_N_829_0\
        );

    \I__8922\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36671\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__36671\,
            I => \Inst_core.Inst_controller.n2717\
        );

    \I__8920\ : CEMux
    port map (
            O => \N__36668\,
            I => \N__36665\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__36665\,
            I => \N__36659\
        );

    \I__8918\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36651\
        );

    \I__8917\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36651\
        );

    \I__8916\ : CascadeMux
    port map (
            O => \N__36662\,
            I => \N__36648\
        );

    \I__8915\ : Span4Mux_h
    port map (
            O => \N__36659\,
            I => \N__36640\
        );

    \I__8914\ : InMux
    port map (
            O => \N__36658\,
            I => \N__36637\
        );

    \I__8913\ : CascadeMux
    port map (
            O => \N__36657\,
            I => \N__36630\
        );

    \I__8912\ : CascadeMux
    port map (
            O => \N__36656\,
            I => \N__36627\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__36651\,
            I => \N__36622\
        );

    \I__8910\ : InMux
    port map (
            O => \N__36648\,
            I => \N__36613\
        );

    \I__8909\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36613\
        );

    \I__8908\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36613\
        );

    \I__8907\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36613\
        );

    \I__8906\ : InMux
    port map (
            O => \N__36644\,
            I => \N__36606\
        );

    \I__8905\ : CEMux
    port map (
            O => \N__36643\,
            I => \N__36603\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__36640\,
            I => \N__36598\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__36637\,
            I => \N__36598\
        );

    \I__8902\ : InMux
    port map (
            O => \N__36636\,
            I => \N__36589\
        );

    \I__8901\ : InMux
    port map (
            O => \N__36635\,
            I => \N__36589\
        );

    \I__8900\ : InMux
    port map (
            O => \N__36634\,
            I => \N__36589\
        );

    \I__8899\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36589\
        );

    \I__8898\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36580\
        );

    \I__8897\ : InMux
    port map (
            O => \N__36627\,
            I => \N__36580\
        );

    \I__8896\ : InMux
    port map (
            O => \N__36626\,
            I => \N__36580\
        );

    \I__8895\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36580\
        );

    \I__8894\ : Span4Mux_s2_v
    port map (
            O => \N__36622\,
            I => \N__36577\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__36613\,
            I => \N__36574\
        );

    \I__8892\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36571\
        );

    \I__8891\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36566\
        );

    \I__8890\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36566\
        );

    \I__8889\ : CEMux
    port map (
            O => \N__36609\,
            I => \N__36558\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__36606\,
            I => \N__36554\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__36603\,
            I => \N__36548\
        );

    \I__8886\ : Span4Mux_h
    port map (
            O => \N__36598\,
            I => \N__36548\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__36589\,
            I => \N__36543\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__36580\,
            I => \N__36543\
        );

    \I__8883\ : Span4Mux_h
    port map (
            O => \N__36577\,
            I => \N__36534\
        );

    \I__8882\ : Span4Mux_s2_v
    port map (
            O => \N__36574\,
            I => \N__36534\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__36571\,
            I => \N__36534\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__36566\,
            I => \N__36534\
        );

    \I__8879\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36525\
        );

    \I__8878\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36525\
        );

    \I__8877\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36525\
        );

    \I__8876\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36525\
        );

    \I__8875\ : CEMux
    port map (
            O => \N__36561\,
            I => \N__36522\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__36558\,
            I => \N__36519\
        );

    \I__8873\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36516\
        );

    \I__8872\ : Span4Mux_v
    port map (
            O => \N__36554\,
            I => \N__36513\
        );

    \I__8871\ : CascadeMux
    port map (
            O => \N__36553\,
            I => \N__36509\
        );

    \I__8870\ : Span4Mux_h
    port map (
            O => \N__36548\,
            I => \N__36503\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__36543\,
            I => \N__36503\
        );

    \I__8868\ : Sp12to4
    port map (
            O => \N__36534\,
            I => \N__36498\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__36525\,
            I => \N__36498\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__36522\,
            I => \N__36495\
        );

    \I__8865\ : Span4Mux_h
    port map (
            O => \N__36519\,
            I => \N__36492\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__36516\,
            I => \N__36489\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__36513\,
            I => \N__36486\
        );

    \I__8862\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36479\
        );

    \I__8861\ : InMux
    port map (
            O => \N__36509\,
            I => \N__36479\
        );

    \I__8860\ : InMux
    port map (
            O => \N__36508\,
            I => \N__36479\
        );

    \I__8859\ : Sp12to4
    port map (
            O => \N__36503\,
            I => \N__36474\
        );

    \I__8858\ : Span12Mux_s1_h
    port map (
            O => \N__36498\,
            I => \N__36474\
        );

    \I__8857\ : Span4Mux_s1_v
    port map (
            O => \N__36495\,
            I => \N__36469\
        );

    \I__8856\ : Span4Mux_v
    port map (
            O => \N__36492\,
            I => \N__36469\
        );

    \I__8855\ : Span4Mux_s1_h
    port map (
            O => \N__36489\,
            I => \N__36462\
        );

    \I__8854\ : Span4Mux_h
    port map (
            O => \N__36486\,
            I => \N__36462\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36462\
        );

    \I__8852\ : Span12Mux_v
    port map (
            O => \N__36474\,
            I => \N__36459\
        );

    \I__8851\ : Odrv4
    port map (
            O => \N__36469\,
            I => \sampleReady\
        );

    \I__8850\ : Odrv4
    port map (
            O => \N__36462\,
            I => \sampleReady\
        );

    \I__8849\ : Odrv12
    port map (
            O => \N__36459\,
            I => \sampleReady\
        );

    \I__8848\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36438\
        );

    \I__8847\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36438\
        );

    \I__8846\ : InMux
    port map (
            O => \N__36450\,
            I => \N__36438\
        );

    \I__8845\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36438\
        );

    \I__8844\ : InMux
    port map (
            O => \N__36448\,
            I => \N__36433\
        );

    \I__8843\ : InMux
    port map (
            O => \N__36447\,
            I => \N__36433\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__36438\,
            I => \Inst_core.n318\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__36433\,
            I => \Inst_core.n318\
        );

    \I__8840\ : CascadeMux
    port map (
            O => \N__36428\,
            I => \Inst_core.Inst_controller.n2717_cascade_\
        );

    \I__8839\ : InMux
    port map (
            O => \N__36425\,
            I => \N__36415\
        );

    \I__8838\ : InMux
    port map (
            O => \N__36424\,
            I => \N__36415\
        );

    \I__8837\ : InMux
    port map (
            O => \N__36423\,
            I => \N__36415\
        );

    \I__8836\ : CascadeMux
    port map (
            O => \N__36422\,
            I => \N__36403\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__36415\,
            I => \N__36396\
        );

    \I__8834\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36393\
        );

    \I__8833\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36390\
        );

    \I__8832\ : InMux
    port map (
            O => \N__36412\,
            I => \N__36375\
        );

    \I__8831\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36375\
        );

    \I__8830\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36375\
        );

    \I__8829\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36375\
        );

    \I__8828\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36375\
        );

    \I__8827\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36375\
        );

    \I__8826\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36375\
        );

    \I__8825\ : InMux
    port map (
            O => \N__36403\,
            I => \N__36370\
        );

    \I__8824\ : InMux
    port map (
            O => \N__36402\,
            I => \N__36370\
        );

    \I__8823\ : InMux
    port map (
            O => \N__36401\,
            I => \N__36363\
        );

    \I__8822\ : InMux
    port map (
            O => \N__36400\,
            I => \N__36363\
        );

    \I__8821\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36363\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__36396\,
            I => \N__36358\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__36393\,
            I => \N__36358\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__36390\,
            I => \N__36353\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__36375\,
            I => \N__36353\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__36370\,
            I => \N__36350\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__36363\,
            I => \N__36347\
        );

    \I__8814\ : Span4Mux_v
    port map (
            O => \N__36358\,
            I => \N__36343\
        );

    \I__8813\ : Span4Mux_s2_v
    port map (
            O => \N__36353\,
            I => \N__36340\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__36350\,
            I => \N__36334\
        );

    \I__8811\ : Span4Mux_v
    port map (
            O => \N__36347\,
            I => \N__36334\
        );

    \I__8810\ : InMux
    port map (
            O => \N__36346\,
            I => \N__36331\
        );

    \I__8809\ : Span4Mux_v
    port map (
            O => \N__36343\,
            I => \N__36326\
        );

    \I__8808\ : Span4Mux_v
    port map (
            O => \N__36340\,
            I => \N__36326\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__36339\,
            I => \N__36322\
        );

    \I__8806\ : Sp12to4
    port map (
            O => \N__36334\,
            I => \N__36310\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__36331\,
            I => \N__36310\
        );

    \I__8804\ : Sp12to4
    port map (
            O => \N__36326\,
            I => \N__36310\
        );

    \I__8803\ : InMux
    port map (
            O => \N__36325\,
            I => \N__36305\
        );

    \I__8802\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36305\
        );

    \I__8801\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36298\
        );

    \I__8800\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36298\
        );

    \I__8799\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36298\
        );

    \I__8798\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36293\
        );

    \I__8797\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36293\
        );

    \I__8796\ : Span12Mux_s11_h
    port map (
            O => \N__36310\,
            I => \N__36290\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__36305\,
            I => send
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__36298\,
            I => send
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__36293\,
            I => send
        );

    \I__8792\ : Odrv12
    port map (
            O => \N__36290\,
            I => send
        );

    \I__8791\ : InMux
    port map (
            O => \N__36281\,
            I => \N__36278\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__36278\,
            I => \Inst_core.Inst_controller.n2\
        );

    \I__8789\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36270\
        );

    \I__8788\ : InMux
    port map (
            O => \N__36274\,
            I => \N__36265\
        );

    \I__8787\ : InMux
    port map (
            O => \N__36273\,
            I => \N__36265\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__36270\,
            I => \Inst_core.Inst_controller.counter_0\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__36265\,
            I => \Inst_core.Inst_controller.counter_0\
        );

    \I__8784\ : InMux
    port map (
            O => \N__36260\,
            I => \bfn_12_12_0_\
        );

    \I__8783\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36252\
        );

    \I__8782\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36249\
        );

    \I__8781\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36246\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__36252\,
            I => \Inst_core.Inst_controller.counter_1\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__36249\,
            I => \Inst_core.Inst_controller.counter_1\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__36246\,
            I => \Inst_core.Inst_controller.counter_1\
        );

    \I__8777\ : InMux
    port map (
            O => \N__36239\,
            I => \Inst_core.Inst_controller.n7845\
        );

    \I__8776\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36231\
        );

    \I__8775\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36228\
        );

    \I__8774\ : InMux
    port map (
            O => \N__36234\,
            I => \N__36225\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__36231\,
            I => \Inst_core.Inst_controller.counter_2\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__36228\,
            I => \Inst_core.Inst_controller.counter_2\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__36225\,
            I => \Inst_core.Inst_controller.counter_2\
        );

    \I__8770\ : InMux
    port map (
            O => \N__36218\,
            I => \Inst_core.Inst_controller.n7846\
        );

    \I__8769\ : CascadeMux
    port map (
            O => \N__36215\,
            I => \N__36212\
        );

    \I__8768\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36208\
        );

    \I__8767\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36205\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__36208\,
            I => \N__36199\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__36205\,
            I => \N__36199\
        );

    \I__8764\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36196\
        );

    \I__8763\ : Span4Mux_h
    port map (
            O => \N__36199\,
            I => \N__36193\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__36196\,
            I => \Inst_core.Inst_controller.counter_3\
        );

    \I__8761\ : Odrv4
    port map (
            O => \N__36193\,
            I => \Inst_core.Inst_controller.counter_3\
        );

    \I__8760\ : InMux
    port map (
            O => \N__36188\,
            I => \Inst_core.Inst_controller.n7847\
        );

    \I__8759\ : InMux
    port map (
            O => \N__36185\,
            I => \N__36181\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__36184\,
            I => \N__36178\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__36181\,
            I => \N__36172\
        );

    \I__8756\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36169\
        );

    \I__8755\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36162\
        );

    \I__8754\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36162\
        );

    \I__8753\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36162\
        );

    \I__8752\ : Span4Mux_v
    port map (
            O => \N__36172\,
            I => \N__36155\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__36169\,
            I => \N__36155\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__36162\,
            I => \N__36152\
        );

    \I__8749\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36147\
        );

    \I__8748\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36147\
        );

    \I__8747\ : Span4Mux_v
    port map (
            O => \N__36155\,
            I => \N__36143\
        );

    \I__8746\ : Span4Mux_v
    port map (
            O => \N__36152\,
            I => \N__36140\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__36147\,
            I => \N__36137\
        );

    \I__8744\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36134\
        );

    \I__8743\ : Odrv4
    port map (
            O => \N__36143\,
            I => cmd_24
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__36140\,
            I => cmd_24
        );

    \I__8741\ : Odrv4
    port map (
            O => \N__36137\,
            I => cmd_24
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__36134\,
            I => cmd_24
        );

    \I__8739\ : CascadeMux
    port map (
            O => \N__36125\,
            I => \N__36122\
        );

    \I__8738\ : InMux
    port map (
            O => \N__36122\,
            I => \N__36119\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__36119\,
            I => \N__36115\
        );

    \I__8736\ : InMux
    port map (
            O => \N__36118\,
            I => \N__36112\
        );

    \I__8735\ : Span4Mux_h
    port map (
            O => \N__36115\,
            I => \N__36109\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__36112\,
            I => \configRegister_16_adj_1344\
        );

    \I__8733\ : Odrv4
    port map (
            O => \N__36109\,
            I => \configRegister_16_adj_1344\
        );

    \I__8732\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36100\
        );

    \I__8731\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36096\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__36100\,
            I => \N__36093\
        );

    \I__8729\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36085\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__36096\,
            I => \N__36080\
        );

    \I__8727\ : Span4Mux_v
    port map (
            O => \N__36093\,
            I => \N__36080\
        );

    \I__8726\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36077\
        );

    \I__8725\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36074\
        );

    \I__8724\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36071\
        );

    \I__8723\ : InMux
    port map (
            O => \N__36089\,
            I => \N__36068\
        );

    \I__8722\ : InMux
    port map (
            O => \N__36088\,
            I => \N__36065\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__36085\,
            I => \N__36062\
        );

    \I__8720\ : Span4Mux_v
    port map (
            O => \N__36080\,
            I => \N__36057\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__36057\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__36074\,
            I => \N__36052\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__36052\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__36068\,
            I => \N__36047\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__36065\,
            I => \N__36047\
        );

    \I__8714\ : Span4Mux_h
    port map (
            O => \N__36062\,
            I => \N__36044\
        );

    \I__8713\ : Span4Mux_s3_h
    port map (
            O => \N__36057\,
            I => \N__36041\
        );

    \I__8712\ : Span4Mux_s3_h
    port map (
            O => \N__36052\,
            I => \N__36038\
        );

    \I__8711\ : Span4Mux_h
    port map (
            O => \N__36047\,
            I => \N__36033\
        );

    \I__8710\ : Span4Mux_h
    port map (
            O => \N__36044\,
            I => \N__36033\
        );

    \I__8709\ : Span4Mux_h
    port map (
            O => \N__36041\,
            I => \N__36030\
        );

    \I__8708\ : Span4Mux_h
    port map (
            O => \N__36038\,
            I => \N__36027\
        );

    \I__8707\ : Odrv4
    port map (
            O => \N__36033\,
            I => wrtrigval_3
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__36030\,
            I => wrtrigval_3
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__36027\,
            I => wrtrigval_3
        );

    \I__8704\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36017\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__36017\,
            I => \N__36014\
        );

    \I__8702\ : Span4Mux_s2_v
    port map (
            O => \N__36014\,
            I => \N__36011\
        );

    \I__8701\ : Span4Mux_v
    port map (
            O => \N__36011\,
            I => \N__36007\
        );

    \I__8700\ : InMux
    port map (
            O => \N__36010\,
            I => \N__36004\
        );

    \I__8699\ : Odrv4
    port map (
            O => \N__36007\,
            I => \valueRegister_0_adj_1376\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__36004\,
            I => \valueRegister_0_adj_1376\
        );

    \I__8697\ : InMux
    port map (
            O => \N__35999\,
            I => \N__35990\
        );

    \I__8696\ : InMux
    port map (
            O => \N__35998\,
            I => \N__35990\
        );

    \I__8695\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35985\
        );

    \I__8694\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35981\
        );

    \I__8693\ : InMux
    port map (
            O => \N__35995\,
            I => \N__35978\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__35990\,
            I => \N__35975\
        );

    \I__8691\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35972\
        );

    \I__8690\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35969\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__35985\,
            I => \N__35966\
        );

    \I__8688\ : InMux
    port map (
            O => \N__35984\,
            I => \N__35963\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__35981\,
            I => \N__35958\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__35978\,
            I => \N__35958\
        );

    \I__8685\ : Span4Mux_s2_v
    port map (
            O => \N__35975\,
            I => \N__35951\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__35972\,
            I => \N__35948\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__35969\,
            I => \N__35945\
        );

    \I__8682\ : Span4Mux_v
    port map (
            O => \N__35966\,
            I => \N__35940\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__35963\,
            I => \N__35940\
        );

    \I__8680\ : Span4Mux_v
    port map (
            O => \N__35958\,
            I => \N__35937\
        );

    \I__8679\ : InMux
    port map (
            O => \N__35957\,
            I => \N__35934\
        );

    \I__8678\ : InMux
    port map (
            O => \N__35956\,
            I => \N__35929\
        );

    \I__8677\ : InMux
    port map (
            O => \N__35955\,
            I => \N__35929\
        );

    \I__8676\ : CascadeMux
    port map (
            O => \N__35954\,
            I => \N__35922\
        );

    \I__8675\ : Span4Mux_v
    port map (
            O => \N__35951\,
            I => \N__35917\
        );

    \I__8674\ : Span4Mux_v
    port map (
            O => \N__35948\,
            I => \N__35917\
        );

    \I__8673\ : Span4Mux_v
    port map (
            O => \N__35945\,
            I => \N__35914\
        );

    \I__8672\ : Span4Mux_v
    port map (
            O => \N__35940\,
            I => \N__35911\
        );

    \I__8671\ : Sp12to4
    port map (
            O => \N__35937\,
            I => \N__35904\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__35934\,
            I => \N__35904\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__35929\,
            I => \N__35904\
        );

    \I__8668\ : InMux
    port map (
            O => \N__35928\,
            I => \N__35901\
        );

    \I__8667\ : InMux
    port map (
            O => \N__35927\,
            I => \N__35896\
        );

    \I__8666\ : InMux
    port map (
            O => \N__35926\,
            I => \N__35896\
        );

    \I__8665\ : InMux
    port map (
            O => \N__35925\,
            I => \N__35893\
        );

    \I__8664\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35890\
        );

    \I__8663\ : Odrv4
    port map (
            O => \N__35917\,
            I => cmd_8
        );

    \I__8662\ : Odrv4
    port map (
            O => \N__35914\,
            I => cmd_8
        );

    \I__8661\ : Odrv4
    port map (
            O => \N__35911\,
            I => cmd_8
        );

    \I__8660\ : Odrv12
    port map (
            O => \N__35904\,
            I => cmd_8
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__35901\,
            I => cmd_8
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__35896\,
            I => cmd_8
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__35893\,
            I => cmd_8
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__35890\,
            I => cmd_8
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__35873\,
            I => \N__35869\
        );

    \I__8654\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35866\
        );

    \I__8653\ : InMux
    port map (
            O => \N__35869\,
            I => \N__35863\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__35866\,
            I => bwd_0
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__35863\,
            I => bwd_0
        );

    \I__8650\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35845\
        );

    \I__8649\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35836\
        );

    \I__8648\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35836\
        );

    \I__8647\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35836\
        );

    \I__8646\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35836\
        );

    \I__8645\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35826\
        );

    \I__8644\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35826\
        );

    \I__8643\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35821\
        );

    \I__8642\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35821\
        );

    \I__8641\ : InMux
    port map (
            O => \N__35849\,
            I => \N__35817\
        );

    \I__8640\ : InMux
    port map (
            O => \N__35848\,
            I => \N__35814\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__35845\,
            I => \N__35808\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__35836\,
            I => \N__35808\
        );

    \I__8637\ : InMux
    port map (
            O => \N__35835\,
            I => \N__35803\
        );

    \I__8636\ : InMux
    port map (
            O => \N__35834\,
            I => \N__35803\
        );

    \I__8635\ : InMux
    port map (
            O => \N__35833\,
            I => \N__35796\
        );

    \I__8634\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35791\
        );

    \I__8633\ : InMux
    port map (
            O => \N__35831\,
            I => \N__35787\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__35826\,
            I => \N__35782\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__35821\,
            I => \N__35782\
        );

    \I__8630\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35779\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__35817\,
            I => \N__35774\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35774\
        );

    \I__8627\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35771\
        );

    \I__8626\ : Span4Mux_v
    port map (
            O => \N__35808\,
            I => \N__35766\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__35803\,
            I => \N__35766\
        );

    \I__8624\ : InMux
    port map (
            O => \N__35802\,
            I => \N__35763\
        );

    \I__8623\ : InMux
    port map (
            O => \N__35801\,
            I => \N__35758\
        );

    \I__8622\ : InMux
    port map (
            O => \N__35800\,
            I => \N__35758\
        );

    \I__8621\ : InMux
    port map (
            O => \N__35799\,
            I => \N__35755\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__35796\,
            I => \N__35752\
        );

    \I__8619\ : InMux
    port map (
            O => \N__35795\,
            I => \N__35749\
        );

    \I__8618\ : InMux
    port map (
            O => \N__35794\,
            I => \N__35746\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__35791\,
            I => \N__35743\
        );

    \I__8616\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35740\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__35787\,
            I => \N__35733\
        );

    \I__8614\ : Span4Mux_v
    port map (
            O => \N__35782\,
            I => \N__35733\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__35779\,
            I => \N__35733\
        );

    \I__8612\ : Span4Mux_v
    port map (
            O => \N__35774\,
            I => \N__35730\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35725\
        );

    \I__8610\ : Span4Mux_v
    port map (
            O => \N__35766\,
            I => \N__35725\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__35763\,
            I => \N__35720\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35720\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35715\
        );

    \I__8606\ : Span4Mux_s3_v
    port map (
            O => \N__35752\,
            I => \N__35715\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__35749\,
            I => \N__35708\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__35746\,
            I => \N__35708\
        );

    \I__8603\ : Span4Mux_v
    port map (
            O => \N__35743\,
            I => \N__35708\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__35740\,
            I => \N__35701\
        );

    \I__8601\ : Span4Mux_v
    port map (
            O => \N__35733\,
            I => \N__35701\
        );

    \I__8600\ : Span4Mux_h
    port map (
            O => \N__35730\,
            I => \N__35701\
        );

    \I__8599\ : Span4Mux_h
    port map (
            O => \N__35725\,
            I => \N__35698\
        );

    \I__8598\ : Span4Mux_s3_v
    port map (
            O => \N__35720\,
            I => \N__35691\
        );

    \I__8597\ : Span4Mux_h
    port map (
            O => \N__35715\,
            I => \N__35691\
        );

    \I__8596\ : Span4Mux_v
    port map (
            O => \N__35708\,
            I => \N__35691\
        );

    \I__8595\ : Span4Mux_h
    port map (
            O => \N__35701\,
            I => \N__35688\
        );

    \I__8594\ : Odrv4
    port map (
            O => \N__35698\,
            I => wrtrigcfg_2
        );

    \I__8593\ : Odrv4
    port map (
            O => \N__35691\,
            I => wrtrigcfg_2
        );

    \I__8592\ : Odrv4
    port map (
            O => \N__35688\,
            I => wrtrigcfg_2
        );

    \I__8591\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35677\
        );

    \I__8590\ : InMux
    port map (
            O => \N__35680\,
            I => \N__35673\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__35677\,
            I => \N__35668\
        );

    \I__8588\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35665\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__35673\,
            I => \N__35662\
        );

    \I__8586\ : InMux
    port map (
            O => \N__35672\,
            I => \N__35659\
        );

    \I__8585\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35656\
        );

    \I__8584\ : Span4Mux_s1_h
    port map (
            O => \N__35668\,
            I => \N__35651\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35651\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__35662\,
            I => \N__35644\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__35659\,
            I => \N__35644\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__35656\,
            I => \N__35644\
        );

    \I__8579\ : Span4Mux_v
    port map (
            O => \N__35651\,
            I => \N__35640\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__35644\,
            I => \N__35637\
        );

    \I__8577\ : InMux
    port map (
            O => \N__35643\,
            I => \N__35634\
        );

    \I__8576\ : Span4Mux_h
    port map (
            O => \N__35640\,
            I => \N__35630\
        );

    \I__8575\ : Span4Mux_h
    port map (
            O => \N__35637\,
            I => \N__35627\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__35634\,
            I => \N__35624\
        );

    \I__8573\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35621\
        );

    \I__8572\ : Odrv4
    port map (
            O => \N__35630\,
            I => cmd_34
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__35627\,
            I => cmd_34
        );

    \I__8570\ : Odrv12
    port map (
            O => \N__35624\,
            I => cmd_34
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__35621\,
            I => cmd_34
        );

    \I__8568\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35607\
        );

    \I__8567\ : CascadeMux
    port map (
            O => \N__35611\,
            I => \N__35602\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__35610\,
            I => \N__35597\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__35607\,
            I => \N__35594\
        );

    \I__8564\ : InMux
    port map (
            O => \N__35606\,
            I => \N__35591\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__35605\,
            I => \N__35588\
        );

    \I__8562\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35585\
        );

    \I__8561\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35582\
        );

    \I__8560\ : CascadeMux
    port map (
            O => \N__35600\,
            I => \N__35579\
        );

    \I__8559\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35575\
        );

    \I__8558\ : Span4Mux_h
    port map (
            O => \N__35594\,
            I => \N__35570\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__35591\,
            I => \N__35570\
        );

    \I__8556\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35567\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__35585\,
            I => \N__35562\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__35582\,
            I => \N__35562\
        );

    \I__8553\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35559\
        );

    \I__8552\ : CascadeMux
    port map (
            O => \N__35578\,
            I => \N__35556\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__35575\,
            I => \N__35553\
        );

    \I__8550\ : Span4Mux_h
    port map (
            O => \N__35570\,
            I => \N__35548\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__35567\,
            I => \N__35548\
        );

    \I__8548\ : Span4Mux_s3_v
    port map (
            O => \N__35562\,
            I => \N__35543\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__35559\,
            I => \N__35543\
        );

    \I__8546\ : InMux
    port map (
            O => \N__35556\,
            I => \N__35540\
        );

    \I__8545\ : Span4Mux_v
    port map (
            O => \N__35553\,
            I => \N__35536\
        );

    \I__8544\ : Span4Mux_s3_v
    port map (
            O => \N__35548\,
            I => \N__35529\
        );

    \I__8543\ : Span4Mux_h
    port map (
            O => \N__35543\,
            I => \N__35529\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__35540\,
            I => \N__35529\
        );

    \I__8541\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35526\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__35536\,
            I => \configRegister_26_adj_1337\
        );

    \I__8539\ : Odrv4
    port map (
            O => \N__35529\,
            I => \configRegister_26_adj_1337\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__35526\,
            I => \configRegister_26_adj_1337\
        );

    \I__8537\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35500\
        );

    \I__8536\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35500\
        );

    \I__8535\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35497\
        );

    \I__8534\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35492\
        );

    \I__8533\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35492\
        );

    \I__8532\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35479\
        );

    \I__8531\ : InMux
    port map (
            O => \N__35513\,
            I => \N__35479\
        );

    \I__8530\ : InMux
    port map (
            O => \N__35512\,
            I => \N__35479\
        );

    \I__8529\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35479\
        );

    \I__8528\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35479\
        );

    \I__8527\ : InMux
    port map (
            O => \N__35509\,
            I => \N__35479\
        );

    \I__8526\ : InMux
    port map (
            O => \N__35508\,
            I => \N__35473\
        );

    \I__8525\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35470\
        );

    \I__8524\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35467\
        );

    \I__8523\ : InMux
    port map (
            O => \N__35505\,
            I => \N__35462\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35453\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__35497\,
            I => \N__35453\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__35492\,
            I => \N__35453\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__35479\,
            I => \N__35453\
        );

    \I__8518\ : InMux
    port map (
            O => \N__35478\,
            I => \N__35448\
        );

    \I__8517\ : InMux
    port map (
            O => \N__35477\,
            I => \N__35448\
        );

    \I__8516\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35445\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__35473\,
            I => \N__35434\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__35470\,
            I => \N__35434\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__35467\,
            I => \N__35434\
        );

    \I__8512\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35427\
        );

    \I__8511\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35427\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__35462\,
            I => \N__35422\
        );

    \I__8509\ : Span4Mux_v
    port map (
            O => \N__35453\,
            I => \N__35422\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__35448\,
            I => \N__35417\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__35445\,
            I => \N__35417\
        );

    \I__8506\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35414\
        );

    \I__8505\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35411\
        );

    \I__8504\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35408\
        );

    \I__8503\ : CascadeMux
    port map (
            O => \N__35441\,
            I => \N__35402\
        );

    \I__8502\ : Span4Mux_v
    port map (
            O => \N__35434\,
            I => \N__35398\
        );

    \I__8501\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35395\
        );

    \I__8500\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35392\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__35427\,
            I => \N__35383\
        );

    \I__8498\ : Span4Mux_s3_h
    port map (
            O => \N__35422\,
            I => \N__35383\
        );

    \I__8497\ : Span4Mux_h
    port map (
            O => \N__35417\,
            I => \N__35383\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__35414\,
            I => \N__35383\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__35411\,
            I => \N__35378\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__35408\,
            I => \N__35378\
        );

    \I__8493\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35375\
        );

    \I__8492\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35366\
        );

    \I__8491\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35366\
        );

    \I__8490\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35366\
        );

    \I__8489\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35366\
        );

    \I__8488\ : Span4Mux_h
    port map (
            O => \N__35398\,
            I => \N__35357\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__35395\,
            I => \N__35357\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__35392\,
            I => \N__35357\
        );

    \I__8485\ : Span4Mux_v
    port map (
            O => \N__35383\,
            I => \N__35354\
        );

    \I__8484\ : Span4Mux_s2_h
    port map (
            O => \N__35378\,
            I => \N__35347\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__35375\,
            I => \N__35347\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35347\
        );

    \I__8481\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35344\
        );

    \I__8480\ : InMux
    port map (
            O => \N__35364\,
            I => \N__35341\
        );

    \I__8479\ : Span4Mux_v
    port map (
            O => \N__35357\,
            I => \N__35338\
        );

    \I__8478\ : Span4Mux_h
    port map (
            O => \N__35354\,
            I => \N__35335\
        );

    \I__8477\ : Span4Mux_h
    port map (
            O => \N__35347\,
            I => \N__35328\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__35344\,
            I => \N__35328\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__35341\,
            I => \N__35328\
        );

    \I__8474\ : Span4Mux_h
    port map (
            O => \N__35338\,
            I => \N__35325\
        );

    \I__8473\ : Span4Mux_h
    port map (
            O => \N__35335\,
            I => \N__35322\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__35328\,
            I => \N__35319\
        );

    \I__8471\ : Odrv4
    port map (
            O => \N__35325\,
            I => wrsize
        );

    \I__8470\ : Odrv4
    port map (
            O => \N__35322\,
            I => wrsize
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__35319\,
            I => wrsize
        );

    \I__8468\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35302\
        );

    \I__8467\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35302\
        );

    \I__8466\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35299\
        );

    \I__8465\ : InMux
    port map (
            O => \N__35309\,
            I => \N__35296\
        );

    \I__8464\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35293\
        );

    \I__8463\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35290\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__35302\,
            I => \N__35286\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__35299\,
            I => \N__35283\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__35296\,
            I => \N__35280\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__35293\,
            I => \N__35277\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__35290\,
            I => \N__35274\
        );

    \I__8457\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35271\
        );

    \I__8456\ : Span4Mux_v
    port map (
            O => \N__35286\,
            I => \N__35267\
        );

    \I__8455\ : Span4Mux_s2_h
    port map (
            O => \N__35283\,
            I => \N__35264\
        );

    \I__8454\ : Span4Mux_s2_h
    port map (
            O => \N__35280\,
            I => \N__35261\
        );

    \I__8453\ : Span4Mux_v
    port map (
            O => \N__35277\,
            I => \N__35254\
        );

    \I__8452\ : Span4Mux_h
    port map (
            O => \N__35274\,
            I => \N__35254\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35254\
        );

    \I__8450\ : InMux
    port map (
            O => \N__35270\,
            I => \N__35251\
        );

    \I__8449\ : Odrv4
    port map (
            O => \N__35267\,
            I => cmd_20
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__35264\,
            I => cmd_20
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__35261\,
            I => cmd_20
        );

    \I__8446\ : Odrv4
    port map (
            O => \N__35254\,
            I => cmd_20
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__35251\,
            I => cmd_20
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__35240\,
            I => \N__35237\
        );

    \I__8443\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35234\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35230\
        );

    \I__8441\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35227\
        );

    \I__8440\ : Span4Mux_v
    port map (
            O => \N__35230\,
            I => \N__35224\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__35227\,
            I => bwd_12
        );

    \I__8438\ : Odrv4
    port map (
            O => \N__35224\,
            I => bwd_12
        );

    \I__8437\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35216\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__35216\,
            I => \N__35212\
        );

    \I__8435\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35209\
        );

    \I__8434\ : Sp12to4
    port map (
            O => \N__35212\,
            I => \N__35204\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__35209\,
            I => \N__35204\
        );

    \I__8432\ : Span12Mux_v
    port map (
            O => \N__35204\,
            I => \N__35201\
        );

    \I__8431\ : Odrv12
    port map (
            O => \N__35201\,
            I => \Inst_core.nstate_1_N_831_0\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__35198\,
            I => \N__35194\
        );

    \I__8429\ : InMux
    port map (
            O => \N__35197\,
            I => \N__35189\
        );

    \I__8428\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35189\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__35189\,
            I => \Inst_core.Inst_controller.n321\
        );

    \I__8426\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35179\
        );

    \I__8425\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35179\
        );

    \I__8424\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35176\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__35179\,
            I => \Inst_core.Inst_controller.nstate_1_N_827_1\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__35176\,
            I => \Inst_core.Inst_controller.nstate_1_N_827_1\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__35171\,
            I => \N__35168\
        );

    \I__8420\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35164\
        );

    \I__8419\ : InMux
    port map (
            O => \N__35167\,
            I => \N__35161\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__35164\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__35161\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8\
        );

    \I__8416\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35152\
        );

    \I__8415\ : InMux
    port map (
            O => \N__35155\,
            I => \N__35149\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__35152\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__35149\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13\
        );

    \I__8412\ : CascadeMux
    port map (
            O => \N__35144\,
            I => \N__35140\
        );

    \I__8411\ : CascadeMux
    port map (
            O => \N__35143\,
            I => \N__35137\
        );

    \I__8410\ : InMux
    port map (
            O => \N__35140\,
            I => \N__35134\
        );

    \I__8409\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35131\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__35134\,
            I => \N__35128\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__35131\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5\
        );

    \I__8406\ : Odrv4
    port map (
            O => \N__35128\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__35123\,
            I => \N__35119\
        );

    \I__8404\ : InMux
    port map (
            O => \N__35122\,
            I => \N__35116\
        );

    \I__8403\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35113\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__35116\,
            I => \N__35110\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__35113\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3\
        );

    \I__8400\ : Odrv4
    port map (
            O => \N__35110\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3\
        );

    \I__8399\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35102\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__35102\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n26\
        );

    \I__8397\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35096\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__35096\,
            I => \N__35092\
        );

    \I__8395\ : InMux
    port map (
            O => \N__35095\,
            I => \N__35089\
        );

    \I__8394\ : Odrv4
    port map (
            O => \N__35092\,
            I => \configRegister_1\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__35089\,
            I => \configRegister_1\
        );

    \I__8392\ : InMux
    port map (
            O => \N__35084\,
            I => \N__35080\
        );

    \I__8391\ : InMux
    port map (
            O => \N__35083\,
            I => \N__35077\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__35080\,
            I => \N__35074\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__35077\,
            I => \configRegister_16\
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__35074\,
            I => \configRegister_16\
        );

    \I__8387\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35064\
        );

    \I__8386\ : InMux
    port map (
            O => \N__35068\,
            I => \N__35061\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__35067\,
            I => \N__35042\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__35064\,
            I => \N__35037\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__35061\,
            I => \N__35037\
        );

    \I__8382\ : InMux
    port map (
            O => \N__35060\,
            I => \N__35034\
        );

    \I__8381\ : InMux
    port map (
            O => \N__35059\,
            I => \N__35031\
        );

    \I__8380\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35026\
        );

    \I__8379\ : InMux
    port map (
            O => \N__35057\,
            I => \N__35026\
        );

    \I__8378\ : InMux
    port map (
            O => \N__35056\,
            I => \N__35023\
        );

    \I__8377\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35018\
        );

    \I__8376\ : InMux
    port map (
            O => \N__35054\,
            I => \N__35018\
        );

    \I__8375\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35014\
        );

    \I__8374\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35011\
        );

    \I__8373\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35006\
        );

    \I__8372\ : InMux
    port map (
            O => \N__35050\,
            I => \N__35006\
        );

    \I__8371\ : InMux
    port map (
            O => \N__35049\,
            I => \N__34997\
        );

    \I__8370\ : InMux
    port map (
            O => \N__35048\,
            I => \N__34997\
        );

    \I__8369\ : InMux
    port map (
            O => \N__35047\,
            I => \N__34997\
        );

    \I__8368\ : InMux
    port map (
            O => \N__35046\,
            I => \N__34997\
        );

    \I__8367\ : InMux
    port map (
            O => \N__35045\,
            I => \N__34992\
        );

    \I__8366\ : InMux
    port map (
            O => \N__35042\,
            I => \N__34989\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__35037\,
            I => \N__34980\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__35034\,
            I => \N__34980\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__34980\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__35026\,
            I => \N__34980\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__35023\,
            I => \N__34977\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__35018\,
            I => \N__34974\
        );

    \I__8359\ : InMux
    port map (
            O => \N__35017\,
            I => \N__34971\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__35014\,
            I => \N__34966\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__35011\,
            I => \N__34966\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__35006\,
            I => \N__34955\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__34997\,
            I => \N__34952\
        );

    \I__8354\ : InMux
    port map (
            O => \N__34996\,
            I => \N__34947\
        );

    \I__8353\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34947\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__34992\,
            I => \N__34944\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__34989\,
            I => \N__34941\
        );

    \I__8350\ : Span4Mux_h
    port map (
            O => \N__34980\,
            I => \N__34936\
        );

    \I__8349\ : Span4Mux_h
    port map (
            O => \N__34977\,
            I => \N__34936\
        );

    \I__8348\ : Span4Mux_h
    port map (
            O => \N__34974\,
            I => \N__34929\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__34971\,
            I => \N__34929\
        );

    \I__8346\ : Span4Mux_h
    port map (
            O => \N__34966\,
            I => \N__34926\
        );

    \I__8345\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34923\
        );

    \I__8344\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34920\
        );

    \I__8343\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34911\
        );

    \I__8342\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34911\
        );

    \I__8341\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34911\
        );

    \I__8340\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34911\
        );

    \I__8339\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34906\
        );

    \I__8338\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34906\
        );

    \I__8337\ : Span4Mux_v
    port map (
            O => \N__34955\,
            I => \N__34901\
        );

    \I__8336\ : Span4Mux_v
    port map (
            O => \N__34952\,
            I => \N__34901\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__34947\,
            I => \N__34898\
        );

    \I__8334\ : Span4Mux_h
    port map (
            O => \N__34944\,
            I => \N__34891\
        );

    \I__8333\ : Span4Mux_h
    port map (
            O => \N__34941\,
            I => \N__34891\
        );

    \I__8332\ : Span4Mux_v
    port map (
            O => \N__34936\,
            I => \N__34891\
        );

    \I__8331\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34886\
        );

    \I__8330\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34886\
        );

    \I__8329\ : Span4Mux_h
    port map (
            O => \N__34929\,
            I => \N__34881\
        );

    \I__8328\ : Span4Mux_h
    port map (
            O => \N__34926\,
            I => \N__34881\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__34923\,
            I => \N__34870\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__34920\,
            I => \N__34870\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__34911\,
            I => \N__34870\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__34906\,
            I => \N__34870\
        );

    \I__8323\ : Sp12to4
    port map (
            O => \N__34901\,
            I => \N__34870\
        );

    \I__8322\ : Span4Mux_v
    port map (
            O => \N__34898\,
            I => \N__34867\
        );

    \I__8321\ : Span4Mux_v
    port map (
            O => \N__34891\,
            I => \N__34864\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__34886\,
            I => \N__34857\
        );

    \I__8319\ : Sp12to4
    port map (
            O => \N__34881\,
            I => \N__34857\
        );

    \I__8318\ : Span12Mux_s8_h
    port map (
            O => \N__34870\,
            I => \N__34857\
        );

    \I__8317\ : Odrv4
    port map (
            O => \N__34867\,
            I => n3753
        );

    \I__8316\ : Odrv4
    port map (
            O => \N__34864\,
            I => n3753
        );

    \I__8315\ : Odrv12
    port map (
            O => \N__34857\,
            I => n3753
        );

    \I__8314\ : CascadeMux
    port map (
            O => \N__34850\,
            I => \N__34847\
        );

    \I__8313\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34836\
        );

    \I__8312\ : InMux
    port map (
            O => \N__34846\,
            I => \N__34827\
        );

    \I__8311\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34827\
        );

    \I__8310\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34827\
        );

    \I__8309\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34827\
        );

    \I__8308\ : CascadeMux
    port map (
            O => \N__34842\,
            I => \N__34822\
        );

    \I__8307\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34814\
        );

    \I__8306\ : CascadeMux
    port map (
            O => \N__34840\,
            I => \N__34811\
        );

    \I__8305\ : CascadeMux
    port map (
            O => \N__34839\,
            I => \N__34806\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__34836\,
            I => \N__34793\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__34827\,
            I => \N__34790\
        );

    \I__8302\ : CascadeMux
    port map (
            O => \N__34826\,
            I => \N__34786\
        );

    \I__8301\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34783\
        );

    \I__8300\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34778\
        );

    \I__8299\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34778\
        );

    \I__8298\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34768\
        );

    \I__8297\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34768\
        );

    \I__8296\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34763\
        );

    \I__8295\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34763\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__34814\,
            I => \N__34760\
        );

    \I__8293\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34757\
        );

    \I__8292\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34754\
        );

    \I__8291\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34747\
        );

    \I__8290\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34747\
        );

    \I__8289\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34747\
        );

    \I__8288\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34744\
        );

    \I__8287\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34739\
        );

    \I__8286\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34739\
        );

    \I__8285\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34736\
        );

    \I__8284\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34733\
        );

    \I__8283\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34730\
        );

    \I__8282\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34725\
        );

    \I__8281\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34725\
        );

    \I__8280\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34722\
        );

    \I__8279\ : Span4Mux_v
    port map (
            O => \N__34793\,
            I => \N__34717\
        );

    \I__8278\ : Span4Mux_v
    port map (
            O => \N__34790\,
            I => \N__34717\
        );

    \I__8277\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34712\
        );

    \I__8276\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34712\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__34783\,
            I => \N__34707\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__34778\,
            I => \N__34707\
        );

    \I__8273\ : CascadeMux
    port map (
            O => \N__34777\,
            I => \N__34703\
        );

    \I__8272\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34695\
        );

    \I__8271\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34692\
        );

    \I__8270\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34687\
        );

    \I__8269\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34687\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34680\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__34763\,
            I => \N__34680\
        );

    \I__8266\ : Span4Mux_h
    port map (
            O => \N__34760\,
            I => \N__34680\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__34757\,
            I => \N__34675\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34675\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__34747\,
            I => \N__34672\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__34744\,
            I => \N__34653\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__34739\,
            I => \N__34653\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__34736\,
            I => \N__34653\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__34733\,
            I => \N__34653\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__34730\,
            I => \N__34653\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__34725\,
            I => \N__34653\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__34722\,
            I => \N__34653\
        );

    \I__8255\ : Span4Mux_h
    port map (
            O => \N__34717\,
            I => \N__34653\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34653\
        );

    \I__8253\ : Span4Mux_s3_h
    port map (
            O => \N__34707\,
            I => \N__34650\
        );

    \I__8252\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34647\
        );

    \I__8251\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34642\
        );

    \I__8250\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34642\
        );

    \I__8249\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34633\
        );

    \I__8248\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34633\
        );

    \I__8247\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34633\
        );

    \I__8246\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34633\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__34695\,
            I => \N__34630\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34627\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__34687\,
            I => \N__34622\
        );

    \I__8242\ : Span4Mux_v
    port map (
            O => \N__34680\,
            I => \N__34622\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__34675\,
            I => \N__34615\
        );

    \I__8240\ : Span4Mux_v
    port map (
            O => \N__34672\,
            I => \N__34615\
        );

    \I__8239\ : Span4Mux_v
    port map (
            O => \N__34653\,
            I => \N__34615\
        );

    \I__8238\ : Span4Mux_v
    port map (
            O => \N__34650\,
            I => \N__34612\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__34647\,
            I => n1
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__34642\,
            I => n1
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__34633\,
            I => n1
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__34630\,
            I => n1
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__34627\,
            I => n1
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__34622\,
            I => n1
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__34615\,
            I => n1
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__34612\,
            I => n1
        );

    \I__8229\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34588\
        );

    \I__8228\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34583\
        );

    \I__8227\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34583\
        );

    \I__8226\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34579\
        );

    \I__8225\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34576\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__34588\,
            I => \N__34573\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__34583\,
            I => \N__34570\
        );

    \I__8222\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34565\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__34579\,
            I => \N__34562\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__34576\,
            I => \N__34555\
        );

    \I__8219\ : Span4Mux_h
    port map (
            O => \N__34573\,
            I => \N__34555\
        );

    \I__8218\ : Span4Mux_s3_v
    port map (
            O => \N__34570\,
            I => \N__34555\
        );

    \I__8217\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34552\
        );

    \I__8216\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34549\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__34565\,
            I => \N__34546\
        );

    \I__8214\ : Span4Mux_h
    port map (
            O => \N__34562\,
            I => \N__34543\
        );

    \I__8213\ : Span4Mux_h
    port map (
            O => \N__34555\,
            I => \N__34540\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__34552\,
            I => cmd_19
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__34549\,
            I => cmd_19
        );

    \I__8210\ : Odrv12
    port map (
            O => \N__34546\,
            I => cmd_19
        );

    \I__8209\ : Odrv4
    port map (
            O => \N__34543\,
            I => cmd_19
        );

    \I__8208\ : Odrv4
    port map (
            O => \N__34540\,
            I => cmd_19
        );

    \I__8207\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34524\
        );

    \I__8206\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34517\
        );

    \I__8205\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34514\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__34524\,
            I => \N__34511\
        );

    \I__8203\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34508\
        );

    \I__8202\ : InMux
    port map (
            O => \N__34522\,
            I => \N__34505\
        );

    \I__8201\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34502\
        );

    \I__8200\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34498\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__34517\,
            I => \N__34495\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__34514\,
            I => \N__34486\
        );

    \I__8197\ : Span4Mux_h
    port map (
            O => \N__34511\,
            I => \N__34486\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__34508\,
            I => \N__34486\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34486\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__34502\,
            I => \N__34483\
        );

    \I__8193\ : CascadeMux
    port map (
            O => \N__34501\,
            I => \N__34480\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__34498\,
            I => \N__34477\
        );

    \I__8191\ : Span4Mux_v
    port map (
            O => \N__34495\,
            I => \N__34474\
        );

    \I__8190\ : Span4Mux_v
    port map (
            O => \N__34486\,
            I => \N__34471\
        );

    \I__8189\ : Span4Mux_s3_h
    port map (
            O => \N__34483\,
            I => \N__34468\
        );

    \I__8188\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34465\
        );

    \I__8187\ : Sp12to4
    port map (
            O => \N__34477\,
            I => \N__34462\
        );

    \I__8186\ : Span4Mux_s1_h
    port map (
            O => \N__34474\,
            I => \N__34459\
        );

    \I__8185\ : Span4Mux_h
    port map (
            O => \N__34471\,
            I => \N__34456\
        );

    \I__8184\ : Span4Mux_h
    port map (
            O => \N__34468\,
            I => \N__34451\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__34465\,
            I => \N__34451\
        );

    \I__8182\ : Span12Mux_s8_h
    port map (
            O => \N__34462\,
            I => \N__34448\
        );

    \I__8181\ : Span4Mux_h
    port map (
            O => \N__34459\,
            I => \N__34443\
        );

    \I__8180\ : Span4Mux_s2_h
    port map (
            O => \N__34456\,
            I => \N__34443\
        );

    \I__8179\ : Span4Mux_v
    port map (
            O => \N__34451\,
            I => \N__34440\
        );

    \I__8178\ : Odrv12
    port map (
            O => \N__34448\,
            I => wrtrigval_1
        );

    \I__8177\ : Odrv4
    port map (
            O => \N__34443\,
            I => wrtrigval_1
        );

    \I__8176\ : Odrv4
    port map (
            O => \N__34440\,
            I => wrtrigval_1
        );

    \I__8175\ : InMux
    port map (
            O => \N__34433\,
            I => \N__34425\
        );

    \I__8174\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34417\
        );

    \I__8173\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34414\
        );

    \I__8172\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34411\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__34429\,
            I => \N__34405\
        );

    \I__8170\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34401\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__34425\,
            I => \N__34398\
        );

    \I__8168\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34395\
        );

    \I__8167\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34392\
        );

    \I__8166\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34389\
        );

    \I__8165\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34386\
        );

    \I__8164\ : InMux
    port map (
            O => \N__34420\,
            I => \N__34383\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__34417\,
            I => \N__34376\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__34414\,
            I => \N__34376\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__34411\,
            I => \N__34376\
        );

    \I__8160\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34373\
        );

    \I__8159\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34368\
        );

    \I__8158\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34368\
        );

    \I__8157\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34363\
        );

    \I__8156\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34363\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__34401\,
            I => \N__34360\
        );

    \I__8154\ : Span4Mux_v
    port map (
            O => \N__34398\,
            I => \N__34357\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__34395\,
            I => \N__34353\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34348\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__34389\,
            I => \N__34348\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__34386\,
            I => \N__34341\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__34383\,
            I => \N__34341\
        );

    \I__8148\ : Span4Mux_v
    port map (
            O => \N__34376\,
            I => \N__34341\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34338\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__34368\,
            I => \N__34335\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__34363\,
            I => \N__34332\
        );

    \I__8144\ : Span4Mux_v
    port map (
            O => \N__34360\,
            I => \N__34327\
        );

    \I__8143\ : Span4Mux_s2_h
    port map (
            O => \N__34357\,
            I => \N__34327\
        );

    \I__8142\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34324\
        );

    \I__8141\ : Span4Mux_v
    port map (
            O => \N__34353\,
            I => \N__34317\
        );

    \I__8140\ : Span4Mux_v
    port map (
            O => \N__34348\,
            I => \N__34317\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__34341\,
            I => \N__34317\
        );

    \I__8138\ : Span4Mux_h
    port map (
            O => \N__34338\,
            I => \N__34308\
        );

    \I__8137\ : Span4Mux_v
    port map (
            O => \N__34335\,
            I => \N__34308\
        );

    \I__8136\ : Span4Mux_v
    port map (
            O => \N__34332\,
            I => \N__34308\
        );

    \I__8135\ : Span4Mux_h
    port map (
            O => \N__34327\,
            I => \N__34308\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__34324\,
            I => cmd_14
        );

    \I__8133\ : Odrv4
    port map (
            O => \N__34317\,
            I => cmd_14
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__34308\,
            I => cmd_14
        );

    \I__8131\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34298\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__34298\,
            I => \N__34295\
        );

    \I__8129\ : Span4Mux_v
    port map (
            O => \N__34295\,
            I => \N__34291\
        );

    \I__8128\ : InMux
    port map (
            O => \N__34294\,
            I => \N__34288\
        );

    \I__8127\ : Odrv4
    port map (
            O => \N__34291\,
            I => \valueRegister_6_adj_1290\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__34288\,
            I => \valueRegister_6_adj_1290\
        );

    \I__8125\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34280\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34276\
        );

    \I__8123\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34273\
        );

    \I__8122\ : Odrv4
    port map (
            O => \N__34276\,
            I => \configRegister_12\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__34273\,
            I => \configRegister_12\
        );

    \I__8120\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34263\
        );

    \I__8119\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34252\
        );

    \I__8118\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34252\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__34263\,
            I => \N__34249\
        );

    \I__8116\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34246\
        );

    \I__8115\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34241\
        );

    \I__8114\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34241\
        );

    \I__8113\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34238\
        );

    \I__8112\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34232\
        );

    \I__8111\ : InMux
    port map (
            O => \N__34257\,
            I => \N__34232\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__34252\,
            I => \N__34228\
        );

    \I__8109\ : Span4Mux_s2_v
    port map (
            O => \N__34249\,
            I => \N__34223\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34216\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__34241\,
            I => \N__34216\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__34238\,
            I => \N__34216\
        );

    \I__8105\ : InMux
    port map (
            O => \N__34237\,
            I => \N__34213\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__34232\,
            I => \N__34210\
        );

    \I__8103\ : InMux
    port map (
            O => \N__34231\,
            I => \N__34207\
        );

    \I__8102\ : Span4Mux_s1_v
    port map (
            O => \N__34228\,
            I => \N__34202\
        );

    \I__8101\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34197\
        );

    \I__8100\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34197\
        );

    \I__8099\ : Span4Mux_v
    port map (
            O => \N__34223\,
            I => \N__34191\
        );

    \I__8098\ : Span4Mux_v
    port map (
            O => \N__34216\,
            I => \N__34191\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__34213\,
            I => \N__34188\
        );

    \I__8096\ : Span4Mux_v
    port map (
            O => \N__34210\,
            I => \N__34183\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__34207\,
            I => \N__34183\
        );

    \I__8094\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34180\
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__34205\,
            I => \N__34176\
        );

    \I__8092\ : Span4Mux_v
    port map (
            O => \N__34202\,
            I => \N__34171\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__34197\,
            I => \N__34171\
        );

    \I__8090\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34168\
        );

    \I__8089\ : Span4Mux_h
    port map (
            O => \N__34191\,
            I => \N__34159\
        );

    \I__8088\ : Span4Mux_v
    port map (
            O => \N__34188\,
            I => \N__34159\
        );

    \I__8087\ : Span4Mux_v
    port map (
            O => \N__34183\,
            I => \N__34159\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__34180\,
            I => \N__34159\
        );

    \I__8085\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34156\
        );

    \I__8084\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34153\
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__34171\,
            I => cmd_9
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__34168\,
            I => cmd_9
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__34159\,
            I => cmd_9
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__34156\,
            I => cmd_9
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__34153\,
            I => cmd_9
        );

    \I__8078\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34139\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__34139\,
            I => \N__34135\
        );

    \I__8076\ : InMux
    port map (
            O => \N__34138\,
            I => \N__34132\
        );

    \I__8075\ : Span4Mux_h
    port map (
            O => \N__34135\,
            I => \N__34129\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__34132\,
            I => bwd_1
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__34129\,
            I => bwd_1
        );

    \I__8072\ : CascadeMux
    port map (
            O => \N__34124\,
            I => \N__34116\
        );

    \I__8071\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34108\
        );

    \I__8070\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34108\
        );

    \I__8069\ : InMux
    port map (
            O => \N__34121\,
            I => \N__34092\
        );

    \I__8068\ : InMux
    port map (
            O => \N__34120\,
            I => \N__34089\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__34119\,
            I => \N__34086\
        );

    \I__8066\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34075\
        );

    \I__8065\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34075\
        );

    \I__8064\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34075\
        );

    \I__8063\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34075\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__34108\,
            I => \N__34072\
        );

    \I__8061\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34067\
        );

    \I__8060\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34067\
        );

    \I__8059\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34064\
        );

    \I__8058\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34057\
        );

    \I__8057\ : InMux
    port map (
            O => \N__34103\,
            I => \N__34057\
        );

    \I__8056\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34057\
        );

    \I__8055\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34050\
        );

    \I__8054\ : InMux
    port map (
            O => \N__34100\,
            I => \N__34050\
        );

    \I__8053\ : InMux
    port map (
            O => \N__34099\,
            I => \N__34050\
        );

    \I__8052\ : CascadeMux
    port map (
            O => \N__34098\,
            I => \N__34047\
        );

    \I__8051\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34041\
        );

    \I__8050\ : InMux
    port map (
            O => \N__34096\,
            I => \N__34041\
        );

    \I__8049\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34038\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34035\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__34089\,
            I => \N__34032\
        );

    \I__8046\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34029\
        );

    \I__8045\ : InMux
    port map (
            O => \N__34085\,
            I => \N__34026\
        );

    \I__8044\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34023\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__34075\,
            I => \N__34020\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__34072\,
            I => \N__34015\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__34067\,
            I => \N__34015\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__34012\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__34057\,
            I => \N__34007\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__34050\,
            I => \N__34007\
        );

    \I__8037\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34002\
        );

    \I__8036\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34002\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__34041\,
            I => \N__33999\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__34038\,
            I => \N__33988\
        );

    \I__8033\ : Span4Mux_h
    port map (
            O => \N__34035\,
            I => \N__33988\
        );

    \I__8032\ : Span4Mux_v
    port map (
            O => \N__34032\,
            I => \N__33988\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__34029\,
            I => \N__33988\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__34026\,
            I => \N__33988\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__34023\,
            I => \N__33985\
        );

    \I__8028\ : Span4Mux_s0_h
    port map (
            O => \N__34020\,
            I => \N__33982\
        );

    \I__8027\ : Span4Mux_v
    port map (
            O => \N__34015\,
            I => \N__33979\
        );

    \I__8026\ : Span4Mux_v
    port map (
            O => \N__34012\,
            I => \N__33974\
        );

    \I__8025\ : Span4Mux_v
    port map (
            O => \N__34007\,
            I => \N__33974\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__34002\,
            I => \N__33971\
        );

    \I__8023\ : Span4Mux_s3_h
    port map (
            O => \N__33999\,
            I => \N__33968\
        );

    \I__8022\ : Span4Mux_v
    port map (
            O => \N__33988\,
            I => \N__33961\
        );

    \I__8021\ : Span4Mux_v
    port map (
            O => \N__33985\,
            I => \N__33961\
        );

    \I__8020\ : Span4Mux_h
    port map (
            O => \N__33982\,
            I => \N__33961\
        );

    \I__8019\ : Span4Mux_v
    port map (
            O => \N__33979\,
            I => \N__33956\
        );

    \I__8018\ : Span4Mux_h
    port map (
            O => \N__33974\,
            I => \N__33956\
        );

    \I__8017\ : Span4Mux_v
    port map (
            O => \N__33971\,
            I => \N__33951\
        );

    \I__8016\ : Span4Mux_h
    port map (
            O => \N__33968\,
            I => \N__33951\
        );

    \I__8015\ : Span4Mux_h
    port map (
            O => \N__33961\,
            I => \N__33948\
        );

    \I__8014\ : Odrv4
    port map (
            O => \N__33956\,
            I => wrtrigcfg_0
        );

    \I__8013\ : Odrv4
    port map (
            O => \N__33951\,
            I => wrtrigcfg_0
        );

    \I__8012\ : Odrv4
    port map (
            O => \N__33948\,
            I => wrtrigcfg_0
        );

    \I__8011\ : CascadeMux
    port map (
            O => \N__33941\,
            I => \N__33937\
        );

    \I__8010\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33932\
        );

    \I__8009\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33929\
        );

    \I__8008\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33923\
        );

    \I__8007\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33923\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__33932\,
            I => \N__33918\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__33929\,
            I => \N__33918\
        );

    \I__8004\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33915\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__33923\,
            I => \N__33908\
        );

    \I__8002\ : Span4Mux_v
    port map (
            O => \N__33918\,
            I => \N__33908\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__33915\,
            I => \N__33905\
        );

    \I__8000\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33902\
        );

    \I__7999\ : InMux
    port map (
            O => \N__33913\,
            I => \N__33899\
        );

    \I__7998\ : Span4Mux_h
    port map (
            O => \N__33908\,
            I => \N__33893\
        );

    \I__7997\ : Span4Mux_v
    port map (
            O => \N__33905\,
            I => \N__33893\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__33902\,
            I => \N__33888\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33888\
        );

    \I__7994\ : InMux
    port map (
            O => \N__33898\,
            I => \N__33885\
        );

    \I__7993\ : Odrv4
    port map (
            O => \N__33893\,
            I => cmd_23
        );

    \I__7992\ : Odrv12
    port map (
            O => \N__33888\,
            I => cmd_23
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__33885\,
            I => cmd_23
        );

    \I__7990\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33875\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__33875\,
            I => \N__33871\
        );

    \I__7988\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33868\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__33871\,
            I => \configRegister_15\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__33868\,
            I => \configRegister_15\
        );

    \I__7985\ : CascadeMux
    port map (
            O => \N__33863\,
            I => \N__33860\
        );

    \I__7984\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33856\
        );

    \I__7983\ : InMux
    port map (
            O => \N__33859\,
            I => \N__33853\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__33856\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__33853\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12\
        );

    \I__7980\ : InMux
    port map (
            O => \N__33848\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7880\
        );

    \I__7979\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33842\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__33842\,
            I => \N__33839\
        );

    \I__7977\ : Span4Mux_s0_h
    port map (
            O => \N__33839\,
            I => \N__33836\
        );

    \I__7976\ : Span4Mux_h
    port map (
            O => \N__33836\,
            I => \N__33832\
        );

    \I__7975\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33829\
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__33832\,
            I => \configRegister_13\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__33829\,
            I => \configRegister_13\
        );

    \I__7972\ : InMux
    port map (
            O => \N__33824\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7881\
        );

    \I__7971\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33818\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__33818\,
            I => \N__33815\
        );

    \I__7969\ : Span4Mux_s0_h
    port map (
            O => \N__33815\,
            I => \N__33811\
        );

    \I__7968\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33808\
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__33811\,
            I => \configRegister_14\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__33808\,
            I => \configRegister_14\
        );

    \I__7965\ : CascadeMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__7964\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33796\
        );

    \I__7963\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33793\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__33796\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__33793\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14\
        );

    \I__7960\ : InMux
    port map (
            O => \N__33788\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7882\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__33785\,
            I => \N__33775\
        );

    \I__7958\ : CascadeMux
    port map (
            O => \N__33784\,
            I => \N__33771\
        );

    \I__7957\ : CascadeMux
    port map (
            O => \N__33783\,
            I => \N__33767\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__33782\,
            I => \N__33762\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__33781\,
            I => \N__33758\
        );

    \I__7954\ : CascadeMux
    port map (
            O => \N__33780\,
            I => \N__33754\
        );

    \I__7953\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33736\
        );

    \I__7952\ : InMux
    port map (
            O => \N__33778\,
            I => \N__33736\
        );

    \I__7951\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33736\
        );

    \I__7950\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33736\
        );

    \I__7949\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33736\
        );

    \I__7948\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33736\
        );

    \I__7947\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33736\
        );

    \I__7946\ : InMux
    port map (
            O => \N__33766\,
            I => \N__33736\
        );

    \I__7945\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33721\
        );

    \I__7944\ : InMux
    port map (
            O => \N__33762\,
            I => \N__33721\
        );

    \I__7943\ : InMux
    port map (
            O => \N__33761\,
            I => \N__33721\
        );

    \I__7942\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33721\
        );

    \I__7941\ : InMux
    port map (
            O => \N__33757\,
            I => \N__33721\
        );

    \I__7940\ : InMux
    port map (
            O => \N__33754\,
            I => \N__33721\
        );

    \I__7939\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33721\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__33736\,
            I => \N__33716\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__33721\,
            I => \N__33716\
        );

    \I__7936\ : Odrv4
    port map (
            O => \N__33716\,
            I => \Inst_core.n1705\
        );

    \I__7935\ : InMux
    port map (
            O => \N__33713\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7883\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__33710\,
            I => \N__33706\
        );

    \I__7933\ : CascadeMux
    port map (
            O => \N__33709\,
            I => \N__33703\
        );

    \I__7932\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33700\
        );

    \I__7931\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33697\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__33700\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__33697\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15\
        );

    \I__7928\ : CEMux
    port map (
            O => \N__33692\,
            I => \N__33688\
        );

    \I__7927\ : CEMux
    port map (
            O => \N__33691\,
            I => \N__33685\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__33688\,
            I => \N__33682\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__33685\,
            I => \N__33679\
        );

    \I__7924\ : Span4Mux_s0_h
    port map (
            O => \N__33682\,
            I => \N__33676\
        );

    \I__7923\ : Span4Mux_s0_h
    port map (
            O => \N__33679\,
            I => \N__33673\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__33676\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4044\
        );

    \I__7921\ : Odrv4
    port map (
            O => \N__33673\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4044\
        );

    \I__7920\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33665\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__33665\,
            I => \N__33661\
        );

    \I__7918\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33658\
        );

    \I__7917\ : Odrv4
    port map (
            O => \N__33661\,
            I => \valueRegister_1_adj_1375\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__33658\,
            I => \valueRegister_1_adj_1375\
        );

    \I__7915\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33648\
        );

    \I__7914\ : CascadeMux
    port map (
            O => \N__33652\,
            I => \N__33642\
        );

    \I__7913\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33639\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__33648\,
            I => \N__33635\
        );

    \I__7911\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33630\
        );

    \I__7910\ : InMux
    port map (
            O => \N__33646\,
            I => \N__33627\
        );

    \I__7909\ : CascadeMux
    port map (
            O => \N__33645\,
            I => \N__33624\
        );

    \I__7908\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33621\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__33639\,
            I => \N__33618\
        );

    \I__7906\ : InMux
    port map (
            O => \N__33638\,
            I => \N__33615\
        );

    \I__7905\ : Span4Mux_v
    port map (
            O => \N__33635\,
            I => \N__33612\
        );

    \I__7904\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33609\
        );

    \I__7903\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33605\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33602\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33599\
        );

    \I__7900\ : InMux
    port map (
            O => \N__33624\,
            I => \N__33596\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__33621\,
            I => \N__33585\
        );

    \I__7898\ : Span4Mux_v
    port map (
            O => \N__33618\,
            I => \N__33585\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__33615\,
            I => \N__33585\
        );

    \I__7896\ : Span4Mux_s3_h
    port map (
            O => \N__33612\,
            I => \N__33585\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__33609\,
            I => \N__33585\
        );

    \I__7894\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33582\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__33605\,
            I => \N__33577\
        );

    \I__7892\ : Span12Mux_s4_h
    port map (
            O => \N__33602\,
            I => \N__33577\
        );

    \I__7891\ : Span12Mux_s11_v
    port map (
            O => \N__33599\,
            I => \N__33574\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33569\
        );

    \I__7889\ : Span4Mux_h
    port map (
            O => \N__33585\,
            I => \N__33569\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__33582\,
            I => \memoryOut_1\
        );

    \I__7887\ : Odrv12
    port map (
            O => \N__33577\,
            I => \memoryOut_1\
        );

    \I__7886\ : Odrv12
    port map (
            O => \N__33574\,
            I => \memoryOut_1\
        );

    \I__7885\ : Odrv4
    port map (
            O => \N__33569\,
            I => \memoryOut_1\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__33560\,
            I => \N__33553\
        );

    \I__7883\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33548\
        );

    \I__7882\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33545\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__33557\,
            I => \N__33542\
        );

    \I__7880\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33539\
        );

    \I__7879\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33535\
        );

    \I__7878\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33532\
        );

    \I__7877\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33529\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__33548\,
            I => \N__33524\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__33545\,
            I => \N__33524\
        );

    \I__7874\ : InMux
    port map (
            O => \N__33542\,
            I => \N__33521\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__33539\,
            I => \N__33518\
        );

    \I__7872\ : InMux
    port map (
            O => \N__33538\,
            I => \N__33515\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__33535\,
            I => \N__33511\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__33532\,
            I => \N__33508\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__33529\,
            I => \N__33505\
        );

    \I__7868\ : Span4Mux_v
    port map (
            O => \N__33524\,
            I => \N__33502\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__33521\,
            I => \N__33495\
        );

    \I__7866\ : Span4Mux_h
    port map (
            O => \N__33518\,
            I => \N__33495\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__33515\,
            I => \N__33495\
        );

    \I__7864\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33492\
        );

    \I__7863\ : Span4Mux_s3_h
    port map (
            O => \N__33511\,
            I => \N__33489\
        );

    \I__7862\ : Span12Mux_s6_v
    port map (
            O => \N__33508\,
            I => \N__33486\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__33505\,
            I => \N__33481\
        );

    \I__7860\ : Span4Mux_h
    port map (
            O => \N__33502\,
            I => \N__33481\
        );

    \I__7859\ : Span4Mux_s2_v
    port map (
            O => \N__33495\,
            I => \N__33478\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__33492\,
            I => \configRegister_26_adj_1377\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__33489\,
            I => \configRegister_26_adj_1377\
        );

    \I__7856\ : Odrv12
    port map (
            O => \N__33486\,
            I => \configRegister_26_adj_1377\
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__33481\,
            I => \configRegister_26_adj_1377\
        );

    \I__7854\ : Odrv4
    port map (
            O => \N__33478\,
            I => \configRegister_26_adj_1377\
        );

    \I__7853\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33464\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__33464\,
            I => \N__33461\
        );

    \I__7851\ : Span4Mux_s0_h
    port map (
            O => \N__33461\,
            I => \N__33458\
        );

    \I__7850\ : Span4Mux_h
    port map (
            O => \N__33458\,
            I => \N__33453\
        );

    \I__7849\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33448\
        );

    \I__7848\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33448\
        );

    \I__7847\ : Odrv4
    port map (
            O => \N__33453\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__33448\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1\
        );

    \I__7845\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33440\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__33440\,
            I => \N__33437\
        );

    \I__7843\ : Span4Mux_s0_h
    port map (
            O => \N__33437\,
            I => \N__33434\
        );

    \I__7842\ : Odrv4
    port map (
            O => \N__33434\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_1\
        );

    \I__7841\ : SRMux
    port map (
            O => \N__33431\,
            I => \N__33428\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__33428\,
            I => \N__33425\
        );

    \I__7839\ : Span4Mux_s1_h
    port map (
            O => \N__33425\,
            I => \N__33422\
        );

    \I__7838\ : Odrv4
    port map (
            O => \N__33422\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4760\
        );

    \I__7837\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33416\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__33416\,
            I => \N__33413\
        );

    \I__7835\ : Span4Mux_v
    port map (
            O => \N__33413\,
            I => \N__33410\
        );

    \I__7834\ : Span4Mux_h
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__7833\ : Odrv4
    port map (
            O => \N__33407\,
            I => \Inst_core.Inst_trigger.stageMatch_2\
        );

    \I__7832\ : InMux
    port map (
            O => \N__33404\,
            I => \N__33401\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__33401\,
            I => \N__33398\
        );

    \I__7830\ : Span4Mux_v
    port map (
            O => \N__33398\,
            I => \N__33395\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__33395\,
            I => \Inst_core.Inst_trigger.stageMatch_3\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__33392\,
            I => \N__33389\
        );

    \I__7827\ : InMux
    port map (
            O => \N__33389\,
            I => \N__33386\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__33386\,
            I => \N__33383\
        );

    \I__7825\ : Span4Mux_v
    port map (
            O => \N__33383\,
            I => \N__33380\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__33380\,
            I => \Inst_core.Inst_trigger.stageMatch_1\
        );

    \I__7823\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33374\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__33374\,
            I => \N__33371\
        );

    \I__7821\ : Odrv12
    port map (
            O => \N__33371\,
            I => \Inst_core.Inst_trigger.stageMatch_0\
        );

    \I__7820\ : CascadeMux
    port map (
            O => \N__33368\,
            I => \N__33365\
        );

    \I__7819\ : InMux
    port map (
            O => \N__33365\,
            I => \N__33359\
        );

    \I__7818\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33359\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__33359\,
            I => \N__33356\
        );

    \I__7816\ : Odrv12
    port map (
            O => \N__33356\,
            I => \Inst_core.Inst_trigger.levelReg_1__N_590\
        );

    \I__7815\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33349\
        );

    \I__7814\ : InMux
    port map (
            O => \N__33352\,
            I => \N__33346\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__33349\,
            I => \N__33343\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__33346\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6\
        );

    \I__7811\ : Odrv12
    port map (
            O => \N__33343\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6\
        );

    \I__7810\ : CascadeMux
    port map (
            O => \N__33338\,
            I => \N__33334\
        );

    \I__7809\ : InMux
    port map (
            O => \N__33337\,
            I => \N__33331\
        );

    \I__7808\ : InMux
    port map (
            O => \N__33334\,
            I => \N__33328\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__33331\,
            I => \N__33325\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__33328\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1\
        );

    \I__7805\ : Odrv4
    port map (
            O => \N__33325\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__33320\,
            I => \N__33317\
        );

    \I__7803\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33313\
        );

    \I__7802\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33310\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33307\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__33310\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4\
        );

    \I__7799\ : Odrv12
    port map (
            O => \N__33307\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4\
        );

    \I__7798\ : CascadeMux
    port map (
            O => \N__33302\,
            I => \N__33298\
        );

    \I__7797\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33295\
        );

    \I__7796\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33292\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__33295\,
            I => \N__33289\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__33292\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0\
        );

    \I__7793\ : Odrv4
    port map (
            O => \N__33289\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0\
        );

    \I__7792\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33281\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__33281\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n28\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__33278\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n25_cascade_\
        );

    \I__7789\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__33272\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n27\
        );

    \I__7787\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33261\
        );

    \I__7786\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33261\
        );

    \I__7785\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33253\
        );

    \I__7784\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33253\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__33261\,
            I => \N__33250\
        );

    \I__7782\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33243\
        );

    \I__7781\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33243\
        );

    \I__7780\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33243\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__33253\,
            I => \N__33240\
        );

    \I__7778\ : Span4Mux_h
    port map (
            O => \N__33250\,
            I => \N__33237\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33234\
        );

    \I__7776\ : Span4Mux_v
    port map (
            O => \N__33240\,
            I => \N__33231\
        );

    \I__7775\ : Odrv4
    port map (
            O => \N__33237\,
            I => \Inst_core.n31_adj_1132\
        );

    \I__7774\ : Odrv12
    port map (
            O => \N__33234\,
            I => \Inst_core.n31_adj_1132\
        );

    \I__7773\ : Odrv4
    port map (
            O => \N__33231\,
            I => \Inst_core.n31_adj_1132\
        );

    \I__7772\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33221\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__33221\,
            I => \N__33217\
        );

    \I__7770\ : InMux
    port map (
            O => \N__33220\,
            I => \N__33214\
        );

    \I__7769\ : Odrv4
    port map (
            O => \N__33217\,
            I => \configRegister_4\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__33214\,
            I => \configRegister_4\
        );

    \I__7767\ : InMux
    port map (
            O => \N__33209\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7872\
        );

    \I__7766\ : InMux
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__33203\,
            I => \N__33199\
        );

    \I__7764\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33196\
        );

    \I__7763\ : Odrv4
    port map (
            O => \N__33199\,
            I => \configRegister_5\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__33196\,
            I => \configRegister_5\
        );

    \I__7761\ : InMux
    port map (
            O => \N__33191\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7873\
        );

    \I__7760\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33185\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__33185\,
            I => \N__33181\
        );

    \I__7758\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33178\
        );

    \I__7757\ : Odrv4
    port map (
            O => \N__33181\,
            I => \configRegister_6\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__33178\,
            I => \configRegister_6\
        );

    \I__7755\ : InMux
    port map (
            O => \N__33173\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7874\
        );

    \I__7754\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33167\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__33167\,
            I => \N__33164\
        );

    \I__7752\ : Span4Mux_v
    port map (
            O => \N__33164\,
            I => \N__33160\
        );

    \I__7751\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33157\
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__33160\,
            I => \configRegister_7\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__33157\,
            I => \configRegister_7\
        );

    \I__7748\ : CascadeMux
    port map (
            O => \N__33152\,
            I => \N__33148\
        );

    \I__7747\ : CascadeMux
    port map (
            O => \N__33151\,
            I => \N__33145\
        );

    \I__7746\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33142\
        );

    \I__7745\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33139\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__33142\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__33139\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7\
        );

    \I__7742\ : InMux
    port map (
            O => \N__33134\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7875\
        );

    \I__7741\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33127\
        );

    \I__7740\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33124\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__33127\,
            I => \N__33121\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__33124\,
            I => \configRegister_8\
        );

    \I__7737\ : Odrv12
    port map (
            O => \N__33121\,
            I => \configRegister_8\
        );

    \I__7736\ : InMux
    port map (
            O => \N__33116\,
            I => \bfn_12_6_0_\
        );

    \I__7735\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33110\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__33110\,
            I => \N__33106\
        );

    \I__7733\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33103\
        );

    \I__7732\ : Odrv4
    port map (
            O => \N__33106\,
            I => \configRegister_9\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__33103\,
            I => \configRegister_9\
        );

    \I__7730\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33094\
        );

    \I__7729\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33091\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__33094\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__33091\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9\
        );

    \I__7726\ : InMux
    port map (
            O => \N__33086\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7877\
        );

    \I__7725\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33080\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__33080\,
            I => \N__33077\
        );

    \I__7723\ : Span4Mux_s3_h
    port map (
            O => \N__33077\,
            I => \N__33073\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33070\
        );

    \I__7721\ : Odrv4
    port map (
            O => \N__33073\,
            I => \configRegister_10\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__33070\,
            I => \configRegister_10\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33058\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33055\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__33058\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__33055\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33050\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7878\
        );

    \I__7713\ : InMux
    port map (
            O => \N__33047\,
            I => \N__33044\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__33044\,
            I => \N__33041\
        );

    \I__7711\ : Span4Mux_v
    port map (
            O => \N__33041\,
            I => \N__33037\
        );

    \I__7710\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33034\
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__33037\,
            I => \configRegister_11\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__33034\,
            I => \configRegister_11\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33029\,
            I => \N__33025\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33028\,
            I => \N__33022\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__33025\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33022\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11\
        );

    \I__7703\ : InMux
    port map (
            O => \N__33017\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7879\
        );

    \I__7702\ : CascadeMux
    port map (
            O => \N__33014\,
            I => \N__33011\
        );

    \I__7701\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33007\
        );

    \I__7700\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33004\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__33007\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__33004\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0\
        );

    \I__7697\ : CascadeMux
    port map (
            O => \N__32999\,
            I => \N__32996\
        );

    \I__7696\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32992\
        );

    \I__7695\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32989\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__32992\,
            I => \N__32986\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__32989\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4\
        );

    \I__7692\ : Odrv4
    port map (
            O => \N__32986\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__32981\,
            I => \N__32978\
        );

    \I__7690\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32974\
        );

    \I__7689\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32971\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__32974\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__32971\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1\
        );

    \I__7686\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32963\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__32963\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n28\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__32960\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n25_cascade_\
        );

    \I__7683\ : InMux
    port map (
            O => \N__32957\,
            I => \N__32954\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__32954\,
            I => \N__32951\
        );

    \I__7681\ : Span4Mux_s3_v
    port map (
            O => \N__32951\,
            I => \N__32944\
        );

    \I__7680\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32935\
        );

    \I__7679\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32935\
        );

    \I__7678\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32935\
        );

    \I__7677\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32935\
        );

    \I__7676\ : Odrv4
    port map (
            O => \N__32944\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n31\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__32935\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n31\
        );

    \I__7674\ : CascadeMux
    port map (
            O => \N__32930\,
            I => \N__32926\
        );

    \I__7673\ : InMux
    port map (
            O => \N__32929\,
            I => \N__32923\
        );

    \I__7672\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32920\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__32923\,
            I => \N__32917\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__32920\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12\
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__32917\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12\
        );

    \I__7668\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32905\
        );

    \I__7666\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32902\
        );

    \I__7665\ : Odrv4
    port map (
            O => \N__32905\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__32902\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2\
        );

    \I__7663\ : CascadeMux
    port map (
            O => \N__32897\,
            I => \N__32893\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__32896\,
            I => \N__32890\
        );

    \I__7661\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32887\
        );

    \I__7660\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32884\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__32887\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__32884\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7\
        );

    \I__7657\ : CascadeMux
    port map (
            O => \N__32879\,
            I => \N__32876\
        );

    \I__7656\ : InMux
    port map (
            O => \N__32876\,
            I => \N__32872\
        );

    \I__7655\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32869\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__32872\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__32869\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10\
        );

    \I__7652\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32861\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__32861\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n27\
        );

    \I__7650\ : CascadeMux
    port map (
            O => \N__32858\,
            I => \N__32855\
        );

    \I__7649\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32851\
        );

    \I__7648\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32848\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__32851\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__32848\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3\
        );

    \I__7645\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32839\
        );

    \I__7644\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32836\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__32839\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__32836\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13\
        );

    \I__7641\ : CascadeMux
    port map (
            O => \N__32831\,
            I => \N__32827\
        );

    \I__7640\ : CascadeMux
    port map (
            O => \N__32830\,
            I => \N__32824\
        );

    \I__7639\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32821\
        );

    \I__7638\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32818\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__32821\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__32818\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__32813\,
            I => \N__32810\
        );

    \I__7634\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32806\
        );

    \I__7633\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32803\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__32806\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__32803\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8\
        );

    \I__7630\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32795\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__32795\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n26\
        );

    \I__7628\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32789\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__32789\,
            I => \N__32785\
        );

    \I__7626\ : InMux
    port map (
            O => \N__32788\,
            I => \N__32782\
        );

    \I__7625\ : Odrv4
    port map (
            O => \N__32785\,
            I => \configRegister_0\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__32782\,
            I => \configRegister_0\
        );

    \I__7623\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32774\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__32774\,
            I => \N__32771\
        );

    \I__7621\ : Span12Mux_s11_v
    port map (
            O => \N__32771\,
            I => \N__32768\
        );

    \I__7620\ : Odrv12
    port map (
            O => \N__32768\,
            I => \Inst_core.n9053\
        );

    \I__7619\ : InMux
    port map (
            O => \N__32765\,
            I => \bfn_12_5_0_\
        );

    \I__7618\ : InMux
    port map (
            O => \N__32762\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7869\
        );

    \I__7617\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32756\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__32756\,
            I => \N__32753\
        );

    \I__7615\ : Span4Mux_v
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__7614\ : Span4Mux_h
    port map (
            O => \N__32750\,
            I => \N__32746\
        );

    \I__7613\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32743\
        );

    \I__7612\ : Odrv4
    port map (
            O => \N__32746\,
            I => \configRegister_2\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__32743\,
            I => \configRegister_2\
        );

    \I__7610\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32734\
        );

    \I__7609\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32731\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__32734\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__32731\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2\
        );

    \I__7606\ : InMux
    port map (
            O => \N__32726\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7870\
        );

    \I__7605\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32720\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__32720\,
            I => \N__32716\
        );

    \I__7603\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32713\
        );

    \I__7602\ : Odrv12
    port map (
            O => \N__32716\,
            I => \configRegister_3\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__32713\,
            I => \configRegister_3\
        );

    \I__7600\ : InMux
    port map (
            O => \N__32708\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7871\
        );

    \I__7599\ : SRMux
    port map (
            O => \N__32705\,
            I => \N__32702\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__32702\,
            I => \N__32699\
        );

    \I__7597\ : Span4Mux_s2_h
    port map (
            O => \N__32699\,
            I => \N__32696\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__32696\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4645\
        );

    \I__7595\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__7593\ : Span4Mux_s1_h
    port map (
            O => \N__32687\,
            I => \N__32684\
        );

    \I__7592\ : Odrv4
    port map (
            O => \N__32684\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_2\
        );

    \I__7591\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32678\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__32678\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_0\
        );

    \I__7589\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32672\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32669\
        );

    \I__7587\ : Span4Mux_h
    port map (
            O => \N__32669\,
            I => \N__32666\
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__32666\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7_adj_1000\
        );

    \I__7585\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32658\
        );

    \I__7584\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32655\
        );

    \I__7583\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32652\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32649\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__32655\,
            I => \Inst_core.Inst_trigger.configRegister_27\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__32652\,
            I => \Inst_core.Inst_trigger.configRegister_27\
        );

    \I__7579\ : Odrv4
    port map (
            O => \N__32649\,
            I => \Inst_core.Inst_trigger.configRegister_27\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__32642\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n8521_cascade_\
        );

    \I__7577\ : CEMux
    port map (
            O => \N__32639\,
            I => \N__32636\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__32636\,
            I => \N__32633\
        );

    \I__7575\ : Span4Mux_s3_v
    port map (
            O => \N__32633\,
            I => \N__32628\
        );

    \I__7574\ : CEMux
    port map (
            O => \N__32632\,
            I => \N__32625\
        );

    \I__7573\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32622\
        );

    \I__7572\ : Span4Mux_s0_h
    port map (
            O => \N__32628\,
            I => \N__32613\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__32625\,
            I => \N__32613\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__32622\,
            I => \N__32613\
        );

    \I__7569\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32610\
        );

    \I__7568\ : CEMux
    port map (
            O => \N__32620\,
            I => \N__32606\
        );

    \I__7567\ : IoSpan4Mux
    port map (
            O => \N__32613\,
            I => \N__32603\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__32610\,
            I => \N__32599\
        );

    \I__7565\ : CEMux
    port map (
            O => \N__32609\,
            I => \N__32596\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__32606\,
            I => \N__32591\
        );

    \I__7563\ : IoSpan4Mux
    port map (
            O => \N__32603\,
            I => \N__32591\
        );

    \I__7562\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32588\
        );

    \I__7561\ : Span4Mux_s3_h
    port map (
            O => \N__32599\,
            I => \N__32585\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32578\
        );

    \I__7559\ : Span4Mux_s3_h
    port map (
            O => \N__32591\,
            I => \N__32578\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__32588\,
            I => \N__32578\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__32585\,
            I => \N__32575\
        );

    \I__7556\ : Span4Mux_h
    port map (
            O => \N__32578\,
            I => \N__32572\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__32575\,
            I => \N__32569\
        );

    \I__7554\ : Span4Mux_v
    port map (
            O => \N__32572\,
            I => \N__32566\
        );

    \I__7553\ : Span4Mux_h
    port map (
            O => \N__32569\,
            I => \N__32563\
        );

    \I__7552\ : Span4Mux_v
    port map (
            O => \N__32566\,
            I => \N__32560\
        );

    \I__7551\ : Odrv4
    port map (
            O => \N__32563\,
            I => \Inst_core.n3670\
        );

    \I__7550\ : Odrv4
    port map (
            O => \N__32560\,
            I => \Inst_core.n3670\
        );

    \I__7549\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32552\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__32552\,
            I => \N__32549\
        );

    \I__7547\ : Span4Mux_s2_v
    port map (
            O => \N__32549\,
            I => \N__32546\
        );

    \I__7546\ : Odrv4
    port map (
            O => \N__32546\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7\
        );

    \I__7545\ : InMux
    port map (
            O => \N__32543\,
            I => \N__32537\
        );

    \I__7544\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32537\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__32537\,
            I => \N__32534\
        );

    \I__7542\ : Span12Mux_s3_h
    port map (
            O => \N__32534\,
            I => \N__32531\
        );

    \I__7541\ : Odrv12
    port map (
            O => \N__32531\,
            I => \Inst_core.Inst_trigger.stageRun_0\
        );

    \I__7540\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32525\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__32525\,
            I => \N__32521\
        );

    \I__7538\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32518\
        );

    \I__7537\ : Span4Mux_s2_h
    port map (
            O => \N__32521\,
            I => \N__32515\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__32518\,
            I => \Inst_core.Inst_trigger.stageRun_3\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__32515\,
            I => \Inst_core.Inst_trigger.stageRun_3\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__32510\,
            I => \N__32507\
        );

    \I__7533\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32500\
        );

    \I__7531\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32497\
        );

    \I__7530\ : Span4Mux_v
    port map (
            O => \N__32500\,
            I => \N__32494\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__32497\,
            I => \Inst_core.stageRun_2\
        );

    \I__7528\ : Odrv4
    port map (
            O => \N__32494\,
            I => \Inst_core.stageRun_2\
        );

    \I__7527\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32485\
        );

    \I__7526\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32482\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__32485\,
            I => \Inst_core.stageRun_1\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__32482\,
            I => \Inst_core.stageRun_1\
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__32477\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n8753_cascade_\
        );

    \I__7522\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32470\
        );

    \I__7521\ : InMux
    port map (
            O => \N__32473\,
            I => \N__32467\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__32470\,
            I => \N__32464\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__32467\,
            I => \N__32461\
        );

    \I__7518\ : Span4Mux_v
    port map (
            O => \N__32464\,
            I => \N__32458\
        );

    \I__7517\ : Span4Mux_v
    port map (
            O => \N__32461\,
            I => \N__32455\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__32458\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n461\
        );

    \I__7515\ : Odrv4
    port map (
            O => \N__32455\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n461\
        );

    \I__7514\ : InMux
    port map (
            O => \N__32450\,
            I => \N__32444\
        );

    \I__7513\ : InMux
    port map (
            O => \N__32449\,
            I => \N__32444\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__32444\,
            I => \N__32441\
        );

    \I__7511\ : Span4Mux_s2_h
    port map (
            O => \N__32441\,
            I => \N__32435\
        );

    \I__7510\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32430\
        );

    \I__7509\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32427\
        );

    \I__7508\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32424\
        );

    \I__7507\ : Span4Mux_v
    port map (
            O => \N__32435\,
            I => \N__32421\
        );

    \I__7506\ : InMux
    port map (
            O => \N__32434\,
            I => \N__32416\
        );

    \I__7505\ : InMux
    port map (
            O => \N__32433\,
            I => \N__32416\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__32430\,
            I => \N__32413\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__32427\,
            I => \N__32408\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__32424\,
            I => \N__32408\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__32421\,
            I => \N__32405\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__32416\,
            I => \Inst_core.state_1\
        );

    \I__7499\ : Odrv12
    port map (
            O => \N__32413\,
            I => \Inst_core.state_1\
        );

    \I__7498\ : Odrv12
    port map (
            O => \N__32408\,
            I => \Inst_core.state_1\
        );

    \I__7497\ : Odrv4
    port map (
            O => \N__32405\,
            I => \Inst_core.state_1\
        );

    \I__7496\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32393\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__32393\,
            I => \N__32389\
        );

    \I__7494\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32386\
        );

    \I__7493\ : Odrv12
    port map (
            O => \N__32389\,
            I => \valueRegister_3_adj_1373\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__32386\,
            I => \valueRegister_3_adj_1373\
        );

    \I__7491\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32378\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__32378\,
            I => \N__32375\
        );

    \I__7489\ : Span12Mux_s4_v
    port map (
            O => \N__32375\,
            I => \N__32370\
        );

    \I__7488\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32365\
        );

    \I__7487\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32365\
        );

    \I__7486\ : Odrv12
    port map (
            O => \N__32370\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__32365\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3\
        );

    \I__7484\ : CascadeMux
    port map (
            O => \N__32360\,
            I => \N__32357\
        );

    \I__7483\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32354\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__32354\,
            I => \N__32348\
        );

    \I__7481\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32345\
        );

    \I__7480\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32340\
        );

    \I__7479\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32334\
        );

    \I__7478\ : Span4Mux_s3_h
    port map (
            O => \N__32348\,
            I => \N__32331\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__32345\,
            I => \N__32328\
        );

    \I__7476\ : InMux
    port map (
            O => \N__32344\,
            I => \N__32323\
        );

    \I__7475\ : InMux
    port map (
            O => \N__32343\,
            I => \N__32323\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__32340\,
            I => \N__32320\
        );

    \I__7473\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32317\
        );

    \I__7472\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32314\
        );

    \I__7471\ : InMux
    port map (
            O => \N__32337\,
            I => \N__32310\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__32334\,
            I => \N__32305\
        );

    \I__7469\ : Span4Mux_v
    port map (
            O => \N__32331\,
            I => \N__32305\
        );

    \I__7468\ : Sp12to4
    port map (
            O => \N__32328\,
            I => \N__32300\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__32323\,
            I => \N__32300\
        );

    \I__7466\ : Span4Mux_s3_v
    port map (
            O => \N__32320\,
            I => \N__32297\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__32317\,
            I => \N__32292\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__32314\,
            I => \N__32292\
        );

    \I__7463\ : InMux
    port map (
            O => \N__32313\,
            I => \N__32289\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__32310\,
            I => \N__32286\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__32305\,
            I => \N__32283\
        );

    \I__7460\ : Span12Mux_s11_v
    port map (
            O => \N__32300\,
            I => \N__32280\
        );

    \I__7459\ : Span4Mux_h
    port map (
            O => \N__32297\,
            I => \N__32275\
        );

    \I__7458\ : Span4Mux_h
    port map (
            O => \N__32292\,
            I => \N__32275\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__32289\,
            I => \memoryOut_3\
        );

    \I__7456\ : Odrv12
    port map (
            O => \N__32286\,
            I => \memoryOut_3\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__32283\,
            I => \memoryOut_3\
        );

    \I__7454\ : Odrv12
    port map (
            O => \N__32280\,
            I => \memoryOut_3\
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__32275\,
            I => \memoryOut_3\
        );

    \I__7452\ : CascadeMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__7451\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32258\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__32258\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_3\
        );

    \I__7449\ : SRMux
    port map (
            O => \N__32255\,
            I => \N__32252\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__32252\,
            I => \N__32249\
        );

    \I__7447\ : Span4Mux_v
    port map (
            O => \N__32249\,
            I => \N__32246\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__32246\,
            I => \N__32243\
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__32243\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4762\
        );

    \I__7444\ : InMux
    port map (
            O => \N__32240\,
            I => \N__32236\
        );

    \I__7443\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32233\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__32236\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__32233\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6\
        );

    \I__7440\ : CEMux
    port map (
            O => \N__32228\,
            I => \N__32225\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__32225\,
            I => \N__32222\
        );

    \I__7438\ : IoSpan4Mux
    port map (
            O => \N__32222\,
            I => \N__32219\
        );

    \I__7437\ : Span4Mux_s0_h
    port map (
            O => \N__32219\,
            I => \N__32216\
        );

    \I__7436\ : Odrv4
    port map (
            O => \N__32216\,
            I => \Inst_core.Inst_sampler.n8687\
        );

    \I__7435\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32210\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__32210\,
            I => \N__32206\
        );

    \I__7433\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32203\
        );

    \I__7432\ : Odrv12
    port map (
            O => \N__32206\,
            I => \valueRegister_0_adj_1336\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__32203\,
            I => \valueRegister_0_adj_1336\
        );

    \I__7430\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32194\
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__32197\,
            I => \N__32191\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__32194\,
            I => \N__32187\
        );

    \I__7427\ : InMux
    port map (
            O => \N__32191\,
            I => \N__32182\
        );

    \I__7426\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32182\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__32187\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__32182\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0\
        );

    \I__7423\ : SRMux
    port map (
            O => \N__32177\,
            I => \N__32174\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__32174\,
            I => \N__32171\
        );

    \I__7421\ : Span4Mux_v
    port map (
            O => \N__32171\,
            I => \N__32168\
        );

    \I__7420\ : Span4Mux_s0_h
    port map (
            O => \N__32168\,
            I => \N__32165\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__32165\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4643\
        );

    \I__7418\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32159\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__32159\,
            I => \N__32156\
        );

    \I__7416\ : Span4Mux_s1_v
    port map (
            O => \N__32156\,
            I => \N__32153\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__32153\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_1\
        );

    \I__7414\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__32147\,
            I => \N__32144\
        );

    \I__7412\ : Odrv12
    port map (
            O => \N__32144\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_2\
        );

    \I__7411\ : CascadeMux
    port map (
            O => \N__32141\,
            I => \N__32138\
        );

    \I__7410\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32135\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__7408\ : Odrv12
    port map (
            O => \N__32132\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_3\
        );

    \I__7407\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32126\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__32126\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_0\
        );

    \I__7405\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32120\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__7403\ : Span4Mux_h
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__7402\ : Span4Mux_v
    port map (
            O => \N__32114\,
            I => \N__32111\
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__32111\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7\
        );

    \I__7400\ : CascadeMux
    port map (
            O => \N__32108\,
            I => \N__32105\
        );

    \I__7399\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32102\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32098\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32094\
        );

    \I__7396\ : Span4Mux_v
    port map (
            O => \N__32098\,
            I => \N__32091\
        );

    \I__7395\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32088\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__32094\,
            I => divider_5
        );

    \I__7393\ : Odrv4
    port map (
            O => \N__32091\,
            I => divider_5
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__32088\,
            I => divider_5
        );

    \I__7391\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32077\
        );

    \I__7390\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32073\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__32077\,
            I => \N__32070\
        );

    \I__7388\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32067\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__32073\,
            I => \N__32060\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__32070\,
            I => \N__32060\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__32067\,
            I => \N__32060\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__32060\,
            I => \Inst_core.Inst_sampler.counter_22\
        );

    \I__7383\ : CascadeMux
    port map (
            O => \N__32057\,
            I => \N__32053\
        );

    \I__7382\ : CascadeMux
    port map (
            O => \N__32056\,
            I => \N__32050\
        );

    \I__7381\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32047\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32043\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32040\
        );

    \I__7378\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32037\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__32032\
        );

    \I__7376\ : Span12Mux_s5_h
    port map (
            O => \N__32040\,
            I => \N__32032\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__32037\,
            I => divider_22
        );

    \I__7374\ : Odrv12
    port map (
            O => \N__32032\,
            I => divider_22
        );

    \I__7373\ : InMux
    port map (
            O => \N__32027\,
            I => \N__32023\
        );

    \I__7372\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32020\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__32023\,
            I => \N__32016\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__32020\,
            I => \N__32013\
        );

    \I__7369\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32010\
        );

    \I__7368\ : Span4Mux_s2_h
    port map (
            O => \N__32016\,
            I => \N__32007\
        );

    \I__7367\ : Span4Mux_s2_h
    port map (
            O => \N__32013\,
            I => \N__32004\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__32010\,
            I => \Inst_core.Inst_sampler.counter_5\
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__32007\,
            I => \Inst_core.Inst_sampler.counter_5\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__32004\,
            I => \Inst_core.Inst_sampler.counter_5\
        );

    \I__7363\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31994\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__31994\,
            I => \Inst_core.Inst_sampler.n34\
        );

    \I__7361\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31988\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31985\
        );

    \I__7359\ : Span4Mux_s3_h
    port map (
            O => \N__31985\,
            I => \N__31982\
        );

    \I__7358\ : Odrv4
    port map (
            O => \N__31982\,
            I => \Inst_core.Inst_sampler.n44\
        );

    \I__7357\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31976\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31973\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__31973\,
            I => \Inst_core.Inst_sampler.n43\
        );

    \I__7354\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31967\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__31967\,
            I => \Inst_core.Inst_sampler.n45\
        );

    \I__7352\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31957\
        );

    \I__7351\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31950\
        );

    \I__7350\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31944\
        );

    \I__7349\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31944\
        );

    \I__7348\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31941\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__31957\,
            I => \N__31938\
        );

    \I__7346\ : IoInMux
    port map (
            O => \N__31956\,
            I => \N__31935\
        );

    \I__7345\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31932\
        );

    \I__7344\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31927\
        );

    \I__7343\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31927\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31924\
        );

    \I__7341\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31921\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__31944\,
            I => \N__31918\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__31941\,
            I => \N__31915\
        );

    \I__7338\ : Span4Mux_v
    port map (
            O => \N__31938\,
            I => \N__31912\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__31935\,
            I => \N__31909\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__31932\,
            I => \N__31904\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__31927\,
            I => \N__31904\
        );

    \I__7334\ : Span4Mux_v
    port map (
            O => \N__31924\,
            I => \N__31897\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__31921\,
            I => \N__31897\
        );

    \I__7332\ : Span4Mux_s2_v
    port map (
            O => \N__31918\,
            I => \N__31897\
        );

    \I__7331\ : Span12Mux_s10_h
    port map (
            O => \N__31915\,
            I => \N__31892\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__31912\,
            I => \N__31889\
        );

    \I__7329\ : Span4Mux_s1_h
    port map (
            O => \N__31909\,
            I => \N__31884\
        );

    \I__7328\ : Span4Mux_h
    port map (
            O => \N__31904\,
            I => \N__31884\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__31897\,
            I => \N__31881\
        );

    \I__7326\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31876\
        );

    \I__7325\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31876\
        );

    \I__7324\ : Span12Mux_v
    port map (
            O => \N__31892\,
            I => \N__31873\
        );

    \I__7323\ : Odrv4
    port map (
            O => \N__31889\,
            I => \ready50_N_581\
        );

    \I__7322\ : Odrv4
    port map (
            O => \N__31884\,
            I => \ready50_N_581\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__31881\,
            I => \ready50_N_581\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__31876\,
            I => \ready50_N_581\
        );

    \I__7319\ : Odrv12
    port map (
            O => \N__31873\,
            I => \ready50_N_581\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__31862\,
            I => \N__31858\
        );

    \I__7317\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31854\
        );

    \I__7316\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31849\
        );

    \I__7315\ : InMux
    port map (
            O => \N__31857\,
            I => \N__31849\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__31854\,
            I => \Inst_core.configRegister_27_adj_1196\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__31849\,
            I => \Inst_core.configRegister_27_adj_1196\
        );

    \I__7312\ : SRMux
    port map (
            O => \N__31844\,
            I => \N__31841\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__31841\,
            I => \N__31838\
        );

    \I__7310\ : Span4Mux_s1_v
    port map (
            O => \N__31838\,
            I => \N__31835\
        );

    \I__7309\ : Odrv4
    port map (
            O => \N__31835\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n8626\
        );

    \I__7308\ : SRMux
    port map (
            O => \N__31832\,
            I => \N__31829\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31826\
        );

    \I__7306\ : Span4Mux_v
    port map (
            O => \N__31826\,
            I => \N__31823\
        );

    \I__7305\ : Span4Mux_v
    port map (
            O => \N__31823\,
            I => \N__31820\
        );

    \I__7304\ : Odrv4
    port map (
            O => \N__31820\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4\
        );

    \I__7303\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31813\
        );

    \I__7302\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31810\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__31813\,
            I => \N__31805\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31805\
        );

    \I__7299\ : Span4Mux_v
    port map (
            O => \N__31805\,
            I => \N__31801\
        );

    \I__7298\ : CascadeMux
    port map (
            O => \N__31804\,
            I => \N__31797\
        );

    \I__7297\ : IoSpan4Mux
    port map (
            O => \N__31801\,
            I => \N__31791\
        );

    \I__7296\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31785\
        );

    \I__7295\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31782\
        );

    \I__7294\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31777\
        );

    \I__7293\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31777\
        );

    \I__7292\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31774\
        );

    \I__7291\ : Span4Mux_s0_h
    port map (
            O => \N__31791\,
            I => \N__31771\
        );

    \I__7290\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31768\
        );

    \I__7289\ : InMux
    port map (
            O => \N__31789\,
            I => \N__31765\
        );

    \I__7288\ : CascadeMux
    port map (
            O => \N__31788\,
            I => \N__31762\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__31785\,
            I => \N__31759\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__31782\,
            I => \N__31756\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__31777\,
            I => \N__31753\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__31774\,
            I => \N__31750\
        );

    \I__7283\ : Span4Mux_h
    port map (
            O => \N__31771\,
            I => \N__31743\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__31768\,
            I => \N__31743\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__31765\,
            I => \N__31743\
        );

    \I__7280\ : InMux
    port map (
            O => \N__31762\,
            I => \N__31740\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__31759\,
            I => \N__31737\
        );

    \I__7278\ : Span12Mux_s4_h
    port map (
            O => \N__31756\,
            I => \N__31734\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__31753\,
            I => \N__31729\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__31750\,
            I => \N__31729\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__31743\,
            I => \N__31726\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__31740\,
            I => \memoryOut_0\
        );

    \I__7273\ : Odrv4
    port map (
            O => \N__31737\,
            I => \memoryOut_0\
        );

    \I__7272\ : Odrv12
    port map (
            O => \N__31734\,
            I => \memoryOut_0\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__31729\,
            I => \memoryOut_0\
        );

    \I__7270\ : Odrv4
    port map (
            O => \N__31726\,
            I => \memoryOut_0\
        );

    \I__7269\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31712\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__31712\,
            I => \N__31709\
        );

    \I__7267\ : Span4Mux_s0_h
    port map (
            O => \N__31709\,
            I => \N__31705\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__31708\,
            I => \N__31702\
        );

    \I__7265\ : Span4Mux_h
    port map (
            O => \N__31705\,
            I => \N__31698\
        );

    \I__7264\ : InMux
    port map (
            O => \N__31702\,
            I => \N__31693\
        );

    \I__7263\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31693\
        );

    \I__7262\ : Odrv4
    port map (
            O => \N__31698\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__31693\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0\
        );

    \I__7260\ : CascadeMux
    port map (
            O => \N__31688\,
            I => \N__31684\
        );

    \I__7259\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31680\
        );

    \I__7258\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31677\
        );

    \I__7257\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31674\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__31680\,
            I => \N__31671\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__31677\,
            I => \N__31668\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__31674\,
            I => \N__31663\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__31671\,
            I => \N__31663\
        );

    \I__7252\ : Span4Mux_s2_h
    port map (
            O => \N__31668\,
            I => \N__31660\
        );

    \I__7251\ : Odrv4
    port map (
            O => \N__31663\,
            I => divider_3
        );

    \I__7250\ : Odrv4
    port map (
            O => \N__31660\,
            I => divider_3
        );

    \I__7249\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31651\
        );

    \I__7248\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31647\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31644\
        );

    \I__7246\ : InMux
    port map (
            O => \N__31650\,
            I => \N__31641\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__31647\,
            I => \N__31634\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__31644\,
            I => \N__31634\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__31641\,
            I => \N__31634\
        );

    \I__7242\ : Odrv4
    port map (
            O => \N__31634\,
            I => \Inst_core.Inst_sampler.counter_6\
        );

    \I__7241\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31628\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__31628\,
            I => \Inst_core.Inst_sampler.n26\
        );

    \I__7239\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__7237\ : Span4Mux_v
    port map (
            O => \N__31619\,
            I => \N__31614\
        );

    \I__7236\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31609\
        );

    \I__7235\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31609\
        );

    \I__7234\ : Odrv4
    port map (
            O => \N__31614\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__31609\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3\
        );

    \I__7232\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31601\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__31601\,
            I => \N__31598\
        );

    \I__7230\ : Span4Mux_s3_h
    port map (
            O => \N__31598\,
            I => \N__31595\
        );

    \I__7229\ : Span4Mux_v
    port map (
            O => \N__31595\,
            I => \N__31591\
        );

    \I__7228\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31588\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__31591\,
            I => \valueRegister_3_adj_1333\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__31588\,
            I => \valueRegister_3_adj_1333\
        );

    \I__7225\ : SRMux
    port map (
            O => \N__31583\,
            I => \N__31580\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__7223\ : Span4Mux_s2_h
    port map (
            O => \N__31577\,
            I => \N__31574\
        );

    \I__7222\ : Span4Mux_s2_v
    port map (
            O => \N__31574\,
            I => \N__31571\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__31571\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4755\
        );

    \I__7220\ : InMux
    port map (
            O => \N__31568\,
            I => \N__31564\
        );

    \I__7219\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31561\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__31564\,
            I => \N__31558\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__31561\,
            I => divider_0
        );

    \I__7216\ : Odrv12
    port map (
            O => \N__31558\,
            I => divider_0
        );

    \I__7215\ : InMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__31550\,
            I => \N__31545\
        );

    \I__7213\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31542\
        );

    \I__7212\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31539\
        );

    \I__7211\ : Span4Mux_s2_h
    port map (
            O => \N__31545\,
            I => \N__31536\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__31542\,
            I => \Inst_core.Inst_sampler.counter_12\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__31539\,
            I => \Inst_core.Inst_sampler.counter_12\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__31536\,
            I => \Inst_core.Inst_sampler.counter_12\
        );

    \I__7207\ : CascadeMux
    port map (
            O => \N__31529\,
            I => \N__31525\
        );

    \I__7206\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31521\
        );

    \I__7205\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31518\
        );

    \I__7204\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31515\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__31521\,
            I => \N__31510\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__31518\,
            I => \N__31510\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__31515\,
            I => divider_12
        );

    \I__7200\ : Odrv12
    port map (
            O => \N__31510\,
            I => divider_12
        );

    \I__7199\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31502\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__31502\,
            I => \N__31499\
        );

    \I__7197\ : Span4Mux_v
    port map (
            O => \N__31499\,
            I => \N__31494\
        );

    \I__7196\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31491\
        );

    \I__7195\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31488\
        );

    \I__7194\ : Span4Mux_s0_h
    port map (
            O => \N__31494\,
            I => \N__31483\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__31491\,
            I => \N__31483\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__31488\,
            I => \Inst_core.Inst_sampler.counter_0\
        );

    \I__7191\ : Odrv4
    port map (
            O => \N__31483\,
            I => \Inst_core.Inst_sampler.counter_0\
        );

    \I__7190\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31475\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__31475\,
            I => \Inst_core.Inst_sampler.n25\
        );

    \I__7188\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31469\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__31469\,
            I => \N__31466\
        );

    \I__7186\ : Span4Mux_h
    port map (
            O => \N__31466\,
            I => \N__31463\
        );

    \I__7185\ : Odrv4
    port map (
            O => \N__31463\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_7\
        );

    \I__7184\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31456\
        );

    \I__7183\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31453\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__31456\,
            I => \N__31450\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__31453\,
            I => \N__31447\
        );

    \I__7180\ : Span4Mux_s3_h
    port map (
            O => \N__31450\,
            I => \N__31444\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__31447\,
            I => \N__31441\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__31444\,
            I => input_c_7
        );

    \I__7177\ : Odrv4
    port map (
            O => \N__31441\,
            I => input_c_7
        );

    \I__7176\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31432\
        );

    \I__7175\ : CascadeMux
    port map (
            O => \N__31435\,
            I => \N__31429\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__31432\,
            I => \N__31425\
        );

    \I__7173\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31422\
        );

    \I__7172\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31419\
        );

    \I__7171\ : Span4Mux_h
    port map (
            O => \N__31425\,
            I => \N__31416\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__31422\,
            I => \N__31413\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__31419\,
            I => \Inst_core.Inst_sync.synchronizedInput_7\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__31416\,
            I => \Inst_core.Inst_sync.synchronizedInput_7\
        );

    \I__7167\ : Odrv12
    port map (
            O => \N__31413\,
            I => \Inst_core.Inst_sync.synchronizedInput_7\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31403\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__31403\,
            I => \N__31399\
        );

    \I__7164\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31394\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__31399\,
            I => \N__31391\
        );

    \I__7162\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31388\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__31397\,
            I => \N__31384\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__31394\,
            I => \N__31380\
        );

    \I__7159\ : Span4Mux_s2_h
    port map (
            O => \N__31391\,
            I => \N__31375\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31375\
        );

    \I__7157\ : InMux
    port map (
            O => \N__31387\,
            I => \N__31371\
        );

    \I__7156\ : InMux
    port map (
            O => \N__31384\,
            I => \N__31365\
        );

    \I__7155\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31361\
        );

    \I__7154\ : Span4Mux_h
    port map (
            O => \N__31380\,
            I => \N__31356\
        );

    \I__7153\ : Span4Mux_v
    port map (
            O => \N__31375\,
            I => \N__31356\
        );

    \I__7152\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31353\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__31371\,
            I => \N__31348\
        );

    \I__7150\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31345\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31342\
        );

    \I__7148\ : InMux
    port map (
            O => \N__31368\,
            I => \N__31339\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__31365\,
            I => \N__31336\
        );

    \I__7146\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31333\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__31361\,
            I => \N__31325\
        );

    \I__7144\ : Span4Mux_h
    port map (
            O => \N__31356\,
            I => \N__31325\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__31353\,
            I => \N__31325\
        );

    \I__7142\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31319\
        );

    \I__7141\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31316\
        );

    \I__7140\ : Span4Mux_v
    port map (
            O => \N__31348\,
            I => \N__31311\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__31345\,
            I => \N__31311\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__31342\,
            I => \N__31306\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31306\
        );

    \I__7136\ : Span4Mux_v
    port map (
            O => \N__31336\,
            I => \N__31303\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__31333\,
            I => \N__31300\
        );

    \I__7134\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31297\
        );

    \I__7133\ : Span4Mux_h
    port map (
            O => \N__31325\,
            I => \N__31294\
        );

    \I__7132\ : CascadeMux
    port map (
            O => \N__31324\,
            I => \N__31291\
        );

    \I__7131\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31288\
        );

    \I__7130\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31285\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__31319\,
            I => \N__31282\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__31316\,
            I => \N__31275\
        );

    \I__7127\ : Span4Mux_v
    port map (
            O => \N__31311\,
            I => \N__31275\
        );

    \I__7126\ : Span4Mux_h
    port map (
            O => \N__31306\,
            I => \N__31275\
        );

    \I__7125\ : Span4Mux_h
    port map (
            O => \N__31303\,
            I => \N__31270\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__31300\,
            I => \N__31270\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31267\
        );

    \I__7122\ : Span4Mux_s1_h
    port map (
            O => \N__31294\,
            I => \N__31264\
        );

    \I__7121\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31261\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31258\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__31285\,
            I => \N__31251\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__31282\,
            I => \N__31251\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__31275\,
            I => \N__31251\
        );

    \I__7116\ : IoSpan4Mux
    port map (
            O => \N__31270\,
            I => \N__31248\
        );

    \I__7115\ : Span4Mux_h
    port map (
            O => \N__31267\,
            I => \N__31243\
        );

    \I__7114\ : Span4Mux_v
    port map (
            O => \N__31264\,
            I => \N__31243\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__31261\,
            I => cmd_13
        );

    \I__7112\ : Odrv12
    port map (
            O => \N__31258\,
            I => cmd_13
        );

    \I__7111\ : Odrv4
    port map (
            O => \N__31251\,
            I => cmd_13
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__31248\,
            I => cmd_13
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__31243\,
            I => cmd_13
        );

    \I__7108\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31229\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__31229\,
            I => \N__31226\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__31226\,
            I => \Inst_core.Inst_sampler.n35\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__31223\,
            I => \N__31220\
        );

    \I__7104\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31217\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31214\
        );

    \I__7102\ : Odrv12
    port map (
            O => \N__31214\,
            I => \Inst_core.Inst_sampler.n36\
        );

    \I__7101\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31208\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31205\
        );

    \I__7099\ : Span4Mux_s2_h
    port map (
            O => \N__31205\,
            I => \N__31202\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__31202\,
            I => \Inst_core.Inst_sampler.n33\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__31199\,
            I => \N__31193\
        );

    \I__7096\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31189\
        );

    \I__7095\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31186\
        );

    \I__7094\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31182\
        );

    \I__7093\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31177\
        );

    \I__7092\ : InMux
    port map (
            O => \N__31192\,
            I => \N__31177\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__31189\,
            I => \N__31172\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__31186\,
            I => \N__31172\
        );

    \I__7089\ : InMux
    port map (
            O => \N__31185\,
            I => \N__31169\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31158\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__31177\,
            I => \N__31158\
        );

    \I__7086\ : Span4Mux_v
    port map (
            O => \N__31172\,
            I => \N__31153\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31169\,
            I => \N__31153\
        );

    \I__7084\ : InMux
    port map (
            O => \N__31168\,
            I => \N__31146\
        );

    \I__7083\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31146\
        );

    \I__7082\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31146\
        );

    \I__7081\ : InMux
    port map (
            O => \N__31165\,
            I => \N__31141\
        );

    \I__7080\ : InMux
    port map (
            O => \N__31164\,
            I => \N__31141\
        );

    \I__7079\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31133\
        );

    \I__7078\ : Span4Mux_v
    port map (
            O => \N__31158\,
            I => \N__31124\
        );

    \I__7077\ : Span4Mux_h
    port map (
            O => \N__31153\,
            I => \N__31124\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__31146\,
            I => \N__31124\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__31141\,
            I => \N__31124\
        );

    \I__7074\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31115\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31139\,
            I => \N__31115\
        );

    \I__7072\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31115\
        );

    \I__7071\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31115\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__31136\,
            I => \N__31107\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__31133\,
            I => \N__31099\
        );

    \I__7068\ : Span4Mux_v
    port map (
            O => \N__31124\,
            I => \N__31094\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__31115\,
            I => \N__31094\
        );

    \I__7066\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31082\
        );

    \I__7065\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31082\
        );

    \I__7064\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31082\
        );

    \I__7063\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31077\
        );

    \I__7062\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31077\
        );

    \I__7061\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31072\
        );

    \I__7060\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31072\
        );

    \I__7059\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31067\
        );

    \I__7058\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31067\
        );

    \I__7057\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31062\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31062\
        );

    \I__7055\ : Span4Mux_v
    port map (
            O => \N__31099\,
            I => \N__31057\
        );

    \I__7054\ : Span4Mux_s3_v
    port map (
            O => \N__31094\,
            I => \N__31057\
        );

    \I__7053\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31054\
        );

    \I__7052\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31051\
        );

    \I__7051\ : InMux
    port map (
            O => \N__31091\,
            I => \N__31048\
        );

    \I__7050\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31043\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31043\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31040\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__31077\,
            I => \N__31035\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__31072\,
            I => \N__31035\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__31067\,
            I => \N__31032\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__31062\,
            I => \N__31028\
        );

    \I__7043\ : Span4Mux_h
    port map (
            O => \N__31057\,
            I => \N__31023\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__31023\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__31051\,
            I => \N__31016\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__31048\,
            I => \N__31016\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__31043\,
            I => \N__31016\
        );

    \I__7038\ : Span4Mux_v
    port map (
            O => \N__31040\,
            I => \N__31013\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__31035\,
            I => \N__31008\
        );

    \I__7036\ : Span4Mux_v
    port map (
            O => \N__31032\,
            I => \N__31008\
        );

    \I__7035\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31005\
        );

    \I__7034\ : Sp12to4
    port map (
            O => \N__31028\,
            I => \N__30998\
        );

    \I__7033\ : Sp12to4
    port map (
            O => \N__31023\,
            I => \N__30998\
        );

    \I__7032\ : Sp12to4
    port map (
            O => \N__31016\,
            I => \N__30998\
        );

    \I__7031\ : Span4Mux_h
    port map (
            O => \N__31013\,
            I => \N__30993\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__31008\,
            I => \N__30993\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__31005\,
            I => \N__30987\
        );

    \I__7028\ : Span12Mux_v
    port map (
            O => \N__30998\,
            I => \N__30987\
        );

    \I__7027\ : Span4Mux_v
    port map (
            O => \N__30993\,
            I => \N__30984\
        );

    \I__7026\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30981\
        );

    \I__7025\ : Odrv12
    port map (
            O => \N__30987\,
            I => \wrDivider\
        );

    \I__7024\ : Odrv4
    port map (
            O => \N__30984\,
            I => \wrDivider\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__30981\,
            I => \wrDivider\
        );

    \I__7022\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30971\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__7020\ : Span4Mux_s2_v
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__30965\,
            I => \Inst_core.Inst_sampler.n8669\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__30962\,
            I => \N__30959\
        );

    \I__7017\ : InMux
    port map (
            O => \N__30959\,
            I => \N__30956\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__30956\,
            I => \N__30953\
        );

    \I__7015\ : Odrv4
    port map (
            O => \N__30953\,
            I => \Inst_core.Inst_sampler.n8671\
        );

    \I__7014\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30947\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__7012\ : Odrv4
    port map (
            O => \N__30944\,
            I => \Inst_core.Inst_sampler.n8673\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__30941\,
            I => \N__30937\
        );

    \I__7010\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30932\
        );

    \I__7009\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30929\
        );

    \I__7008\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30925\
        );

    \I__7007\ : InMux
    port map (
            O => \N__30935\,
            I => \N__30918\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__30932\,
            I => \N__30913\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__30929\,
            I => \N__30913\
        );

    \I__7004\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30910\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30906\
        );

    \I__7002\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30903\
        );

    \I__7001\ : InMux
    port map (
            O => \N__30923\,
            I => \N__30900\
        );

    \I__7000\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30895\
        );

    \I__6999\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30895\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__30918\,
            I => \N__30892\
        );

    \I__6997\ : Span4Mux_v
    port map (
            O => \N__30913\,
            I => \N__30889\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__30910\,
            I => \N__30886\
        );

    \I__6995\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30883\
        );

    \I__6994\ : Span4Mux_v
    port map (
            O => \N__30906\,
            I => \N__30880\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__30903\,
            I => \N__30875\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__30900\,
            I => \N__30875\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__30895\,
            I => \N__30872\
        );

    \I__6990\ : Span4Mux_v
    port map (
            O => \N__30892\,
            I => \N__30867\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__30889\,
            I => \N__30867\
        );

    \I__6988\ : Span12Mux_v
    port map (
            O => \N__30886\,
            I => \N__30864\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__30883\,
            I => \N__30859\
        );

    \I__6986\ : Span4Mux_v
    port map (
            O => \N__30880\,
            I => \N__30859\
        );

    \I__6985\ : Span4Mux_v
    port map (
            O => \N__30875\,
            I => \N__30854\
        );

    \I__6984\ : Span4Mux_h
    port map (
            O => \N__30872\,
            I => \N__30854\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__30867\,
            I => \memoryOut_2\
        );

    \I__6982\ : Odrv12
    port map (
            O => \N__30864\,
            I => \memoryOut_2\
        );

    \I__6981\ : Odrv4
    port map (
            O => \N__30859\,
            I => \memoryOut_2\
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__30854\,
            I => \memoryOut_2\
        );

    \I__6979\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30842\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__30842\,
            I => \N__30839\
        );

    \I__6977\ : Span4Mux_s2_h
    port map (
            O => \N__30839\,
            I => \N__30835\
        );

    \I__6976\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30832\
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__30835\,
            I => \valueRegister_2_adj_1334\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__30832\,
            I => \valueRegister_2_adj_1334\
        );

    \I__6973\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30824\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__30824\,
            I => \N__30820\
        );

    \I__6971\ : CascadeMux
    port map (
            O => \N__30823\,
            I => \N__30817\
        );

    \I__6970\ : Span4Mux_h
    port map (
            O => \N__30820\,
            I => \N__30813\
        );

    \I__6969\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30808\
        );

    \I__6968\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30808\
        );

    \I__6967\ : Odrv4
    port map (
            O => \N__30813\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__30808\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2\
        );

    \I__6965\ : SRMux
    port map (
            O => \N__30803\,
            I => \N__30800\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__30800\,
            I => \N__30797\
        );

    \I__6963\ : Span4Mux_v
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__6962\ : Span4Mux_h
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__6961\ : Span4Mux_v
    port map (
            O => \N__30791\,
            I => \N__30788\
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__30788\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4754\
        );

    \I__6959\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30781\
        );

    \I__6958\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30778\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__30781\,
            I => \N__30775\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30772\
        );

    \I__6955\ : Span4Mux_h
    port map (
            O => \N__30775\,
            I => \N__30768\
        );

    \I__6954\ : Span4Mux_v
    port map (
            O => \N__30772\,
            I => \N__30765\
        );

    \I__6953\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30762\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__30768\,
            I => \N__30759\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__30765\,
            I => \N__30756\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__30762\,
            I => divider_11
        );

    \I__6949\ : Odrv4
    port map (
            O => \N__30759\,
            I => divider_11
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__30756\,
            I => divider_11
        );

    \I__6947\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30746\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30742\
        );

    \I__6945\ : InMux
    port map (
            O => \N__30745\,
            I => \N__30739\
        );

    \I__6944\ : Span4Mux_s2_h
    port map (
            O => \N__30742\,
            I => \N__30736\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__30739\,
            I => \Inst_core.Inst_sampler.counter_23\
        );

    \I__6942\ : Odrv4
    port map (
            O => \N__30736\,
            I => \Inst_core.Inst_sampler.counter_23\
        );

    \I__6941\ : CascadeMux
    port map (
            O => \N__30731\,
            I => \N__30728\
        );

    \I__6940\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30722\
        );

    \I__6939\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30722\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__30722\,
            I => \N__30718\
        );

    \I__6937\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30715\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__30718\,
            I => \N__30712\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__30715\,
            I => \Inst_core.Inst_sampler.counter_11\
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__30712\,
            I => \Inst_core.Inst_sampler.counter_11\
        );

    \I__6933\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30704\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__30704\,
            I => \N__30700\
        );

    \I__6931\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30696\
        );

    \I__6930\ : Span4Mux_s2_h
    port map (
            O => \N__30700\,
            I => \N__30693\
        );

    \I__6929\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30690\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__30696\,
            I => \Inst_core.Inst_sampler.counter_2\
        );

    \I__6927\ : Odrv4
    port map (
            O => \N__30693\,
            I => \Inst_core.Inst_sampler.counter_2\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__30690\,
            I => \Inst_core.Inst_sampler.counter_2\
        );

    \I__6925\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30680\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__30680\,
            I => \N__30677\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__30677\,
            I => \Inst_core.Inst_sampler.n8606\
        );

    \I__6922\ : CascadeMux
    port map (
            O => \N__30674\,
            I => \Inst_core.Inst_sampler.n3_cascade_\
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__30671\,
            I => \N__30667\
        );

    \I__6920\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30661\
        );

    \I__6919\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30661\
        );

    \I__6918\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30658\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__30661\,
            I => \N__30655\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__30658\,
            I => divider_23
        );

    \I__6915\ : Odrv12
    port map (
            O => \N__30655\,
            I => divider_23
        );

    \I__6914\ : InMux
    port map (
            O => \N__30650\,
            I => \N__30647\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__6912\ : Odrv4
    port map (
            O => \N__30644\,
            I => \Inst_core.Inst_sampler.n8618\
        );

    \I__6911\ : CascadeMux
    port map (
            O => \N__30641\,
            I => \Inst_core.Inst_sampler.n8656_cascade_\
        );

    \I__6910\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30633\
        );

    \I__6909\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30630\
        );

    \I__6908\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30627\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__30633\,
            I => \N__30622\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__30630\,
            I => \N__30622\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__30627\,
            I => divider_1
        );

    \I__6904\ : Odrv12
    port map (
            O => \N__30622\,
            I => divider_1
        );

    \I__6903\ : InMux
    port map (
            O => \N__30617\,
            I => \N__30613\
        );

    \I__6902\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30610\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__30613\,
            I => \N__30606\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__30610\,
            I => \N__30603\
        );

    \I__6899\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30600\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__30606\,
            I => \N__30595\
        );

    \I__6897\ : Span4Mux_v
    port map (
            O => \N__30603\,
            I => \N__30595\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__30600\,
            I => \Inst_core.Inst_sampler.counter_18\
        );

    \I__6895\ : Odrv4
    port map (
            O => \N__30595\,
            I => \Inst_core.Inst_sampler.counter_18\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__30590\,
            I => \N__30587\
        );

    \I__6893\ : InMux
    port map (
            O => \N__30587\,
            I => \N__30584\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__30584\,
            I => \N__30580\
        );

    \I__6891\ : InMux
    port map (
            O => \N__30583\,
            I => \N__30576\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__30580\,
            I => \N__30573\
        );

    \I__6889\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30570\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__30576\,
            I => \N__30567\
        );

    \I__6887\ : Span4Mux_s0_h
    port map (
            O => \N__30573\,
            I => \N__30564\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__30570\,
            I => divider_18
        );

    \I__6885\ : Odrv4
    port map (
            O => \N__30567\,
            I => divider_18
        );

    \I__6884\ : Odrv4
    port map (
            O => \N__30564\,
            I => divider_18
        );

    \I__6883\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30552\
        );

    \I__6882\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30549\
        );

    \I__6881\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30546\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__30552\,
            I => \N__30541\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30541\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__30546\,
            I => \Inst_core.Inst_sampler.counter_1\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__30541\,
            I => \Inst_core.Inst_sampler.counter_1\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30533\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__30533\,
            I => \N__30530\
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__30530\,
            I => \Inst_core.Inst_sampler.n28\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__30527\,
            I => \Inst_core.Inst_sampler.n27_cascade_\
        );

    \I__6872\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30519\
        );

    \I__6871\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30516\
        );

    \I__6870\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30513\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30508\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30508\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__30513\,
            I => divider_6
        );

    \I__6866\ : Odrv12
    port map (
            O => \N__30508\,
            I => divider_6
        );

    \I__6865\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30498\
        );

    \I__6864\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30495\
        );

    \I__6863\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30492\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__30498\,
            I => \N__30487\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30487\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__30492\,
            I => \Inst_core.Inst_sampler.counter_3\
        );

    \I__6859\ : Odrv4
    port map (
            O => \N__30487\,
            I => \Inst_core.Inst_sampler.counter_3\
        );

    \I__6858\ : SRMux
    port map (
            O => \N__30482\,
            I => \N__30479\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__30479\,
            I => \N__30476\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__30476\,
            I => \N__30473\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__30473\,
            I => \N__30470\
        );

    \I__6854\ : Odrv4
    port map (
            O => \N__30470\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4747\
        );

    \I__6853\ : CascadeMux
    port map (
            O => \N__30467\,
            I => \N__30463\
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__30466\,
            I => \N__30458\
        );

    \I__6851\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30453\
        );

    \I__6850\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30449\
        );

    \I__6849\ : InMux
    port map (
            O => \N__30461\,
            I => \N__30446\
        );

    \I__6848\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30443\
        );

    \I__6847\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30439\
        );

    \I__6846\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30436\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__30453\,
            I => \N__30433\
        );

    \I__6844\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30429\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__30449\,
            I => \N__30426\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__30446\,
            I => \N__30423\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__30443\,
            I => \N__30420\
        );

    \I__6840\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30417\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__30439\,
            I => \N__30414\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30409\
        );

    \I__6837\ : Span4Mux_h
    port map (
            O => \N__30433\,
            I => \N__30409\
        );

    \I__6836\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30406\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__30429\,
            I => \N__30402\
        );

    \I__6834\ : Span4Mux_v
    port map (
            O => \N__30426\,
            I => \N__30397\
        );

    \I__6833\ : Span4Mux_s3_v
    port map (
            O => \N__30423\,
            I => \N__30397\
        );

    \I__6832\ : Span4Mux_h
    port map (
            O => \N__30420\,
            I => \N__30394\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__30417\,
            I => \N__30391\
        );

    \I__6830\ : Sp12to4
    port map (
            O => \N__30414\,
            I => \N__30386\
        );

    \I__6829\ : Sp12to4
    port map (
            O => \N__30409\,
            I => \N__30386\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__30406\,
            I => \N__30383\
        );

    \I__6827\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30380\
        );

    \I__6826\ : Span4Mux_h
    port map (
            O => \N__30402\,
            I => \N__30373\
        );

    \I__6825\ : Span4Mux_h
    port map (
            O => \N__30397\,
            I => \N__30373\
        );

    \I__6824\ : Span4Mux_v
    port map (
            O => \N__30394\,
            I => \N__30373\
        );

    \I__6823\ : Span12Mux_s5_h
    port map (
            O => \N__30391\,
            I => \N__30366\
        );

    \I__6822\ : Span12Mux_s11_v
    port map (
            O => \N__30386\,
            I => \N__30366\
        );

    \I__6821\ : Span12Mux_s6_h
    port map (
            O => \N__30383\,
            I => \N__30366\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__30380\,
            I => \memoryOut_6\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__30373\,
            I => \memoryOut_6\
        );

    \I__6818\ : Odrv12
    port map (
            O => \N__30366\,
            I => \memoryOut_6\
        );

    \I__6817\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30354\
        );

    \I__6816\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30351\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__30357\,
            I => \N__30348\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__30354\,
            I => \N__30339\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__30351\,
            I => \N__30339\
        );

    \I__6812\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30336\
        );

    \I__6811\ : CascadeMux
    port map (
            O => \N__30347\,
            I => \N__30333\
        );

    \I__6810\ : CascadeMux
    port map (
            O => \N__30346\,
            I => \N__30329\
        );

    \I__6809\ : InMux
    port map (
            O => \N__30345\,
            I => \N__30326\
        );

    \I__6808\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30323\
        );

    \I__6807\ : Span4Mux_h
    port map (
            O => \N__30339\,
            I => \N__30320\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__30336\,
            I => \N__30317\
        );

    \I__6805\ : InMux
    port map (
            O => \N__30333\,
            I => \N__30314\
        );

    \I__6804\ : InMux
    port map (
            O => \N__30332\,
            I => \N__30311\
        );

    \I__6803\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30308\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__30326\,
            I => \N__30305\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__30323\,
            I => \N__30302\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__30320\,
            I => \N__30297\
        );

    \I__6799\ : Span4Mux_h
    port map (
            O => \N__30317\,
            I => \N__30297\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__30314\,
            I => \N__30293\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__30311\,
            I => \N__30288\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__30308\,
            I => \N__30288\
        );

    \I__6795\ : Span4Mux_s2_v
    port map (
            O => \N__30305\,
            I => \N__30285\
        );

    \I__6794\ : Span4Mux_s2_h
    port map (
            O => \N__30302\,
            I => \N__30282\
        );

    \I__6793\ : Span4Mux_v
    port map (
            O => \N__30297\,
            I => \N__30279\
        );

    \I__6792\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30276\
        );

    \I__6791\ : Span4Mux_v
    port map (
            O => \N__30293\,
            I => \N__30273\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__30288\,
            I => \N__30268\
        );

    \I__6789\ : Span4Mux_v
    port map (
            O => \N__30285\,
            I => \N__30268\
        );

    \I__6788\ : Span4Mux_v
    port map (
            O => \N__30282\,
            I => \N__30263\
        );

    \I__6787\ : Span4Mux_h
    port map (
            O => \N__30279\,
            I => \N__30263\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__30276\,
            I => \configRegister_26_adj_1297\
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__30273\,
            I => \configRegister_26_adj_1297\
        );

    \I__6784\ : Odrv4
    port map (
            O => \N__30268\,
            I => \configRegister_26_adj_1297\
        );

    \I__6783\ : Odrv4
    port map (
            O => \N__30263\,
            I => \configRegister_26_adj_1297\
        );

    \I__6782\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__30251\,
            I => \N__30248\
        );

    \I__6780\ : Span4Mux_s2_h
    port map (
            O => \N__30248\,
            I => \N__30245\
        );

    \I__6779\ : Span4Mux_h
    port map (
            O => \N__30245\,
            I => \N__30241\
        );

    \I__6778\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30238\
        );

    \I__6777\ : Odrv4
    port map (
            O => \N__30241\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__30238\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6\
        );

    \I__6775\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30230\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__30230\,
            I => \N__30227\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__30227\,
            I => \N__30224\
        );

    \I__6772\ : Odrv4
    port map (
            O => \N__30224\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_6\
        );

    \I__6771\ : SRMux
    port map (
            O => \N__30221\,
            I => \N__30218\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__30218\,
            I => \N__30215\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__30215\,
            I => \N__30212\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__30212\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4751\
        );

    \I__6767\ : InMux
    port map (
            O => \N__30209\,
            I => \N__30206\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__30206\,
            I => \N__30202\
        );

    \I__6765\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30199\
        );

    \I__6764\ : Span4Mux_v
    port map (
            O => \N__30202\,
            I => \N__30196\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__30199\,
            I => fwd_0
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__30196\,
            I => fwd_0
        );

    \I__6761\ : CascadeMux
    port map (
            O => \N__30191\,
            I => \N__30188\
        );

    \I__6760\ : InMux
    port map (
            O => \N__30188\,
            I => \N__30184\
        );

    \I__6759\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30181\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__30184\,
            I => \N__30178\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__30181\,
            I => fwd_2
        );

    \I__6756\ : Odrv12
    port map (
            O => \N__30178\,
            I => fwd_2
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__30173\,
            I => \N__30170\
        );

    \I__6754\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__6752\ : Span4Mux_v
    port map (
            O => \N__30164\,
            I => \N__30161\
        );

    \I__6751\ : Span4Mux_h
    port map (
            O => \N__30161\,
            I => \N__30158\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__30158\,
            I => \Inst_core.Inst_controller.n16\
        );

    \I__6749\ : IoInMux
    port map (
            O => \N__30155\,
            I => \N__30151\
        );

    \I__6748\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30148\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__30151\,
            I => \N__30145\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__30148\,
            I => \N__30141\
        );

    \I__6745\ : Span4Mux_s1_h
    port map (
            O => \N__30145\,
            I => \N__30138\
        );

    \I__6744\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30135\
        );

    \I__6743\ : Span12Mux_s10_h
    port map (
            O => \N__30141\,
            I => \N__30132\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__30138\,
            I => debugleds_c_1
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__30135\,
            I => debugleds_c_1
        );

    \I__6740\ : Odrv12
    port map (
            O => \N__30132\,
            I => debugleds_c_1
        );

    \I__6739\ : CascadeMux
    port map (
            O => \N__30125\,
            I => \Inst_core.n4_cascade_\
        );

    \I__6738\ : CascadeMux
    port map (
            O => \N__30122\,
            I => \Inst_core.Inst_controller.n3907_cascade_\
        );

    \I__6737\ : CascadeMux
    port map (
            O => \N__30119\,
            I => \N__30116\
        );

    \I__6736\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30110\
        );

    \I__6735\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30107\
        );

    \I__6734\ : InMux
    port map (
            O => \N__30114\,
            I => \N__30104\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__30113\,
            I => \N__30101\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__30110\,
            I => \N__30095\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30095\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__30104\,
            I => \N__30092\
        );

    \I__6729\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30089\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30100\,
            I => \N__30086\
        );

    \I__6727\ : Span4Mux_h
    port map (
            O => \N__30095\,
            I => \N__30082\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__30092\,
            I => \N__30079\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30089\,
            I => \N__30076\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__30086\,
            I => \N__30073\
        );

    \I__6723\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30070\
        );

    \I__6722\ : Span4Mux_v
    port map (
            O => \N__30082\,
            I => \N__30065\
        );

    \I__6721\ : Span4Mux_v
    port map (
            O => \N__30079\,
            I => \N__30062\
        );

    \I__6720\ : Span4Mux_v
    port map (
            O => \N__30076\,
            I => \N__30059\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__30073\,
            I => \N__30054\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__30070\,
            I => \N__30054\
        );

    \I__6717\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30051\
        );

    \I__6716\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30048\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__30065\,
            I => cmd_22
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__30062\,
            I => cmd_22
        );

    \I__6713\ : Odrv4
    port map (
            O => \N__30059\,
            I => cmd_22
        );

    \I__6712\ : Odrv4
    port map (
            O => \N__30054\,
            I => cmd_22
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__30051\,
            I => cmd_22
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__30048\,
            I => cmd_22
        );

    \I__6709\ : InMux
    port map (
            O => \N__30035\,
            I => \N__30030\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__30034\,
            I => \N__30027\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__30033\,
            I => \N__30024\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__30030\,
            I => \N__30020\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30017\
        );

    \I__6704\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30012\
        );

    \I__6703\ : InMux
    port map (
            O => \N__30023\,
            I => \N__30012\
        );

    \I__6702\ : Span4Mux_v
    port map (
            O => \N__30020\,
            I => \N__30009\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__30017\,
            I => cmd_26
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__30012\,
            I => cmd_26
        );

    \I__6699\ : Odrv4
    port map (
            O => \N__30009\,
            I => cmd_26
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__30002\,
            I => \N__29998\
        );

    \I__6697\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29993\
        );

    \I__6696\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29993\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__29993\,
            I => \N__29990\
        );

    \I__6694\ : Span4Mux_s2_h
    port map (
            O => \N__29990\,
            I => \N__29985\
        );

    \I__6693\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29980\
        );

    \I__6692\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29980\
        );

    \I__6691\ : Odrv4
    port map (
            O => \N__29985\,
            I => cmd_27
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__29980\,
            I => cmd_27
        );

    \I__6689\ : CascadeMux
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__6688\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29968\
        );

    \I__6687\ : CascadeMux
    port map (
            O => \N__29971\,
            I => \N__29965\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__29968\,
            I => \N__29962\
        );

    \I__6685\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29959\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__29962\,
            I => \N__29955\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__29959\,
            I => \N__29952\
        );

    \I__6682\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29949\
        );

    \I__6681\ : Span4Mux_v
    port map (
            O => \N__29955\,
            I => \N__29946\
        );

    \I__6680\ : Span4Mux_h
    port map (
            O => \N__29952\,
            I => \N__29943\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__29949\,
            I => divider_19
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__29946\,
            I => divider_19
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__29943\,
            I => divider_19
        );

    \I__6676\ : InMux
    port map (
            O => \N__29936\,
            I => \N__29933\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__29933\,
            I => \N__29929\
        );

    \I__6674\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29926\
        );

    \I__6673\ : Span4Mux_s3_h
    port map (
            O => \N__29929\,
            I => \N__29923\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__29926\,
            I => bwd_2
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__29923\,
            I => bwd_2
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__29918\,
            I => \N__29915\
        );

    \I__6669\ : InMux
    port map (
            O => \N__29915\,
            I => \N__29911\
        );

    \I__6668\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29908\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__29911\,
            I => \N__29905\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__29908\,
            I => bwd_13
        );

    \I__6665\ : Odrv12
    port map (
            O => \N__29905\,
            I => bwd_13
        );

    \I__6664\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29897\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__29897\,
            I => \N__29894\
        );

    \I__6662\ : Span4Mux_s3_h
    port map (
            O => \N__29894\,
            I => \N__29891\
        );

    \I__6661\ : Odrv4
    port map (
            O => \N__29891\,
            I => \Inst_core.Inst_controller.n18_adj_990\
        );

    \I__6660\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29885\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__29885\,
            I => \N__29882\
        );

    \I__6658\ : Odrv12
    port map (
            O => \N__29882\,
            I => \Inst_core.Inst_controller.n20\
        );

    \I__6657\ : CascadeMux
    port map (
            O => \N__29879\,
            I => \Inst_core.Inst_controller.n17_cascade_\
        );

    \I__6656\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29873\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__29873\,
            I => \N__29870\
        );

    \I__6654\ : Span4Mux_s2_h
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__6653\ : Odrv4
    port map (
            O => \N__29867\,
            I => \Inst_core.Inst_controller.n30\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__29864\,
            I => \Inst_core.Inst_controller.n29_cascade_\
        );

    \I__6651\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29858\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__29858\,
            I => \N__29855\
        );

    \I__6649\ : Span4Mux_h
    port map (
            O => \N__29855\,
            I => \N__29852\
        );

    \I__6648\ : Odrv4
    port map (
            O => \N__29852\,
            I => \Inst_core.Inst_controller.n6693\
        );

    \I__6647\ : InMux
    port map (
            O => \N__29849\,
            I => \N__29845\
        );

    \I__6646\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29842\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__29845\,
            I => \N__29839\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__29842\,
            I => \Inst_core.Inst_controller.bwd_14\
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__29839\,
            I => \Inst_core.Inst_controller.bwd_14\
        );

    \I__6642\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__29831\,
            I => \Inst_core.Inst_controller.n19\
        );

    \I__6640\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__29825\,
            I => \N__29821\
        );

    \I__6638\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29818\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__29821\,
            I => \valueRegister_2_adj_1294\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__29818\,
            I => \valueRegister_2_adj_1294\
        );

    \I__6635\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29810\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__29810\,
            I => \N__29806\
        );

    \I__6633\ : CascadeMux
    port map (
            O => \N__29809\,
            I => \N__29803\
        );

    \I__6632\ : Span4Mux_s2_h
    port map (
            O => \N__29806\,
            I => \N__29799\
        );

    \I__6631\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29794\
        );

    \I__6630\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29794\
        );

    \I__6629\ : Odrv4
    port map (
            O => \N__29799\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__29794\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2\
        );

    \I__6627\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29786\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__29786\,
            I => \N__29783\
        );

    \I__6625\ : Odrv12
    port map (
            O => \N__29783\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_2\
        );

    \I__6624\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29776\
        );

    \I__6623\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29773\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__29776\,
            I => \N__29770\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__29773\,
            I => \maskRegister_6_adj_1282\
        );

    \I__6620\ : Odrv12
    port map (
            O => \N__29770\,
            I => \maskRegister_6_adj_1282\
        );

    \I__6619\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29759\
        );

    \I__6618\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29759\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__29759\,
            I => \N__29753\
        );

    \I__6616\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29746\
        );

    \I__6615\ : InMux
    port map (
            O => \N__29757\,
            I => \N__29746\
        );

    \I__6614\ : CascadeMux
    port map (
            O => \N__29756\,
            I => \N__29742\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__29753\,
            I => \N__29739\
        );

    \I__6612\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29736\
        );

    \I__6611\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29733\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__29746\,
            I => \N__29730\
        );

    \I__6609\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29725\
        );

    \I__6608\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29725\
        );

    \I__6607\ : Odrv4
    port map (
            O => \N__29739\,
            I => cmd_31
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__29736\,
            I => cmd_31
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__29733\,
            I => cmd_31
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__29730\,
            I => cmd_31
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__29725\,
            I => cmd_31
        );

    \I__6602\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29708\
        );

    \I__6601\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29699\
        );

    \I__6600\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29699\
        );

    \I__6599\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29699\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__29708\,
            I => \N__29696\
        );

    \I__6597\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29693\
        );

    \I__6596\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29688\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__29699\,
            I => \N__29685\
        );

    \I__6594\ : Span4Mux_h
    port map (
            O => \N__29696\,
            I => \N__29680\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29680\
        );

    \I__6592\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29672\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__29691\,
            I => \N__29668\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__29688\,
            I => \N__29665\
        );

    \I__6589\ : Span4Mux_v
    port map (
            O => \N__29685\,
            I => \N__29662\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__29680\,
            I => \N__29659\
        );

    \I__6587\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29656\
        );

    \I__6586\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29653\
        );

    \I__6585\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29650\
        );

    \I__6584\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29647\
        );

    \I__6583\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29644\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__29672\,
            I => \N__29641\
        );

    \I__6581\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29638\
        );

    \I__6580\ : InMux
    port map (
            O => \N__29668\,
            I => \N__29635\
        );

    \I__6579\ : Span4Mux_v
    port map (
            O => \N__29665\,
            I => \N__29626\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__29662\,
            I => \N__29626\
        );

    \I__6577\ : Span4Mux_s2_v
    port map (
            O => \N__29659\,
            I => \N__29626\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__29656\,
            I => \N__29626\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__29653\,
            I => \N__29616\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__29650\,
            I => \N__29616\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__29647\,
            I => \N__29616\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__29644\,
            I => \N__29611\
        );

    \I__6571\ : Span4Mux_v
    port map (
            O => \N__29641\,
            I => \N__29611\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__29638\,
            I => \N__29606\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__29635\,
            I => \N__29606\
        );

    \I__6568\ : Sp12to4
    port map (
            O => \N__29626\,
            I => \N__29603\
        );

    \I__6567\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29598\
        );

    \I__6566\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29598\
        );

    \I__6565\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29595\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__29616\,
            I => \N__29592\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__29611\,
            I => \N__29589\
        );

    \I__6562\ : Span12Mux_s6_h
    port map (
            O => \N__29606\,
            I => \N__29584\
        );

    \I__6561\ : Span12Mux_s7_v
    port map (
            O => \N__29603\,
            I => \N__29584\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__29598\,
            I => cmd_10
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__29595\,
            I => cmd_10
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__29592\,
            I => cmd_10
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__29589\,
            I => cmd_10
        );

    \I__6556\ : Odrv12
    port map (
            O => \N__29584\,
            I => cmd_10
        );

    \I__6555\ : CascadeMux
    port map (
            O => \N__29573\,
            I => \N__29570\
        );

    \I__6554\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__29567\,
            I => \N__29563\
        );

    \I__6552\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29560\
        );

    \I__6551\ : Odrv12
    port map (
            O => \N__29563\,
            I => \valueRegister_2_adj_1374\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__29560\,
            I => \valueRegister_2_adj_1374\
        );

    \I__6549\ : InMux
    port map (
            O => \N__29555\,
            I => \N__29549\
        );

    \I__6548\ : InMux
    port map (
            O => \N__29554\,
            I => \N__29549\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__29549\,
            I => \N__29545\
        );

    \I__6546\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29542\
        );

    \I__6545\ : Span4Mux_h
    port map (
            O => \N__29545\,
            I => \N__29535\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__29542\,
            I => \N__29535\
        );

    \I__6543\ : InMux
    port map (
            O => \N__29541\,
            I => \N__29532\
        );

    \I__6542\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29529\
        );

    \I__6541\ : Span4Mux_s3_h
    port map (
            O => \N__29535\,
            I => \N__29520\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__29532\,
            I => \N__29520\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__29529\,
            I => \N__29520\
        );

    \I__6538\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29517\
        );

    \I__6537\ : CascadeMux
    port map (
            O => \N__29527\,
            I => \N__29514\
        );

    \I__6536\ : Span4Mux_v
    port map (
            O => \N__29520\,
            I => \N__29510\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__29517\,
            I => \N__29507\
        );

    \I__6534\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29502\
        );

    \I__6533\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29502\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__29510\,
            I => cmd_25
        );

    \I__6531\ : Odrv12
    port map (
            O => \N__29507\,
            I => cmd_25
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__29502\,
            I => cmd_25
        );

    \I__6529\ : CascadeMux
    port map (
            O => \N__29495\,
            I => \N__29491\
        );

    \I__6528\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29484\
        );

    \I__6527\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29484\
        );

    \I__6526\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29479\
        );

    \I__6525\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29476\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29472\
        );

    \I__6523\ : InMux
    port map (
            O => \N__29483\,
            I => \N__29467\
        );

    \I__6522\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29467\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__29479\,
            I => \N__29464\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__29476\,
            I => \N__29461\
        );

    \I__6519\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29458\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__29472\,
            I => \N__29452\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__29467\,
            I => \N__29452\
        );

    \I__6516\ : Span4Mux_v
    port map (
            O => \N__29464\,
            I => \N__29449\
        );

    \I__6515\ : Span4Mux_s2_h
    port map (
            O => \N__29461\,
            I => \N__29444\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__29458\,
            I => \N__29444\
        );

    \I__6513\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29441\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__29452\,
            I => \N__29438\
        );

    \I__6511\ : Span4Mux_v
    port map (
            O => \N__29449\,
            I => \N__29433\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__29444\,
            I => \N__29433\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__29441\,
            I => \N__29430\
        );

    \I__6508\ : Span4Mux_v
    port map (
            O => \N__29438\,
            I => \N__29427\
        );

    \I__6507\ : Span4Mux_h
    port map (
            O => \N__29433\,
            I => \N__29424\
        );

    \I__6506\ : Span4Mux_h
    port map (
            O => \N__29430\,
            I => \N__29421\
        );

    \I__6505\ : Odrv4
    port map (
            O => \N__29427\,
            I => wrtrigval_2
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__29424\,
            I => wrtrigval_2
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__29421\,
            I => wrtrigval_2
        );

    \I__6502\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29410\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29407\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__29410\,
            I => \N__29404\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__29407\,
            I => \configRegister_17\
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__29404\,
            I => \configRegister_17\
        );

    \I__6497\ : CascadeMux
    port map (
            O => \N__29399\,
            I => \N__29396\
        );

    \I__6496\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29391\
        );

    \I__6495\ : InMux
    port map (
            O => \N__29395\,
            I => \N__29388\
        );

    \I__6494\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29385\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__29391\,
            I => \N__29379\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__29388\,
            I => \N__29374\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__29385\,
            I => \N__29374\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29369\
        );

    \I__6489\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29369\
        );

    \I__6488\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29366\
        );

    \I__6487\ : Span4Mux_h
    port map (
            O => \N__29379\,
            I => \N__29363\
        );

    \I__6486\ : Span4Mux_h
    port map (
            O => \N__29374\,
            I => \N__29356\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__29369\,
            I => \N__29356\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29356\
        );

    \I__6483\ : Span4Mux_v
    port map (
            O => \N__29363\,
            I => \N__29351\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__29356\,
            I => \N__29348\
        );

    \I__6481\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29345\
        );

    \I__6480\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29342\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__29351\,
            I => cmd_21
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__29348\,
            I => cmd_21
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__29345\,
            I => cmd_21
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__29342\,
            I => cmd_21
        );

    \I__6475\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29327\
        );

    \I__6474\ : InMux
    port map (
            O => \N__29332\,
            I => \N__29321\
        );

    \I__6473\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29315\
        );

    \I__6472\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29312\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__29327\,
            I => \N__29307\
        );

    \I__6470\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29304\
        );

    \I__6469\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29301\
        );

    \I__6468\ : CascadeMux
    port map (
            O => \N__29324\,
            I => \N__29296\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__29321\,
            I => \N__29287\
        );

    \I__6466\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29284\
        );

    \I__6465\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29279\
        );

    \I__6464\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29279\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__29315\,
            I => \N__29274\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__29312\,
            I => \N__29274\
        );

    \I__6461\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29271\
        );

    \I__6460\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29268\
        );

    \I__6459\ : Span4Mux_v
    port map (
            O => \N__29307\,
            I => \N__29262\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__29304\,
            I => \N__29262\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__29301\,
            I => \N__29259\
        );

    \I__6456\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29254\
        );

    \I__6455\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29254\
        );

    \I__6454\ : InMux
    port map (
            O => \N__29296\,
            I => \N__29243\
        );

    \I__6453\ : InMux
    port map (
            O => \N__29295\,
            I => \N__29243\
        );

    \I__6452\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29243\
        );

    \I__6451\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29240\
        );

    \I__6450\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29237\
        );

    \I__6449\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29234\
        );

    \I__6448\ : InMux
    port map (
            O => \N__29290\,
            I => \N__29231\
        );

    \I__6447\ : Span4Mux_h
    port map (
            O => \N__29287\,
            I => \N__29224\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__29284\,
            I => \N__29224\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29224\
        );

    \I__6444\ : Span4Mux_h
    port map (
            O => \N__29274\,
            I => \N__29217\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29217\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__29268\,
            I => \N__29217\
        );

    \I__6441\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29214\
        );

    \I__6440\ : Span4Mux_v
    port map (
            O => \N__29262\,
            I => \N__29211\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__29259\,
            I => \N__29206\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__29254\,
            I => \N__29206\
        );

    \I__6437\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29197\
        );

    \I__6436\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29197\
        );

    \I__6435\ : InMux
    port map (
            O => \N__29251\,
            I => \N__29197\
        );

    \I__6434\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29197\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__29243\,
            I => \N__29194\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29240\,
            I => \N__29187\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__29237\,
            I => \N__29187\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__29234\,
            I => \N__29187\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29184\
        );

    \I__6428\ : Span4Mux_v
    port map (
            O => \N__29224\,
            I => \N__29179\
        );

    \I__6427\ : Span4Mux_v
    port map (
            O => \N__29217\,
            I => \N__29179\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29176\
        );

    \I__6425\ : Span4Mux_h
    port map (
            O => \N__29211\,
            I => \N__29171\
        );

    \I__6424\ : Span4Mux_h
    port map (
            O => \N__29206\,
            I => \N__29171\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29164\
        );

    \I__6422\ : Span4Mux_s3_v
    port map (
            O => \N__29194\,
            I => \N__29164\
        );

    \I__6421\ : Span4Mux_v
    port map (
            O => \N__29187\,
            I => \N__29164\
        );

    \I__6420\ : Span4Mux_v
    port map (
            O => \N__29184\,
            I => \N__29159\
        );

    \I__6419\ : Span4Mux_h
    port map (
            O => \N__29179\,
            I => \N__29159\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__29176\,
            I => \N__29152\
        );

    \I__6417\ : Span4Mux_v
    port map (
            O => \N__29171\,
            I => \N__29152\
        );

    \I__6416\ : Span4Mux_h
    port map (
            O => \N__29164\,
            I => \N__29152\
        );

    \I__6415\ : Odrv4
    port map (
            O => \N__29159\,
            I => wrtrigcfg_1
        );

    \I__6414\ : Odrv4
    port map (
            O => \N__29152\,
            I => wrtrigcfg_1
        );

    \I__6413\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__29144\,
            I => \N__29140\
        );

    \I__6411\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29137\
        );

    \I__6410\ : Odrv12
    port map (
            O => \N__29140\,
            I => \configRegister_14_adj_1306\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__29137\,
            I => \configRegister_14_adj_1306\
        );

    \I__6408\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29124\
        );

    \I__6407\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29119\
        );

    \I__6406\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29116\
        );

    \I__6405\ : InMux
    port map (
            O => \N__29129\,
            I => \N__29111\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__29128\,
            I => \N__29104\
        );

    \I__6403\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29101\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__29124\,
            I => \N__29098\
        );

    \I__6401\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29092\
        );

    \I__6400\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29092\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__29119\,
            I => \N__29089\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__29116\,
            I => \N__29086\
        );

    \I__6397\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29083\
        );

    \I__6396\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29080\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__29111\,
            I => \N__29077\
        );

    \I__6394\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29074\
        );

    \I__6393\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29071\
        );

    \I__6392\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29068\
        );

    \I__6391\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29065\
        );

    \I__6390\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29060\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__29101\,
            I => \N__29057\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__29098\,
            I => \N__29054\
        );

    \I__6387\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29051\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__29092\,
            I => \N__29044\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__29089\,
            I => \N__29044\
        );

    \I__6384\ : Span4Mux_v
    port map (
            O => \N__29086\,
            I => \N__29044\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__29083\,
            I => \N__29041\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29036\
        );

    \I__6381\ : Span4Mux_v
    port map (
            O => \N__29077\,
            I => \N__29036\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__29074\,
            I => \N__29027\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29027\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29027\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29027\
        );

    \I__6376\ : InMux
    port map (
            O => \N__29064\,
            I => \N__29024\
        );

    \I__6375\ : InMux
    port map (
            O => \N__29063\,
            I => \N__29021\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__29060\,
            I => \N__29018\
        );

    \I__6373\ : Span4Mux_h
    port map (
            O => \N__29057\,
            I => \N__29015\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__29054\,
            I => \N__29012\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__29051\,
            I => \N__29007\
        );

    \I__6370\ : Span4Mux_h
    port map (
            O => \N__29044\,
            I => \N__29007\
        );

    \I__6369\ : Span4Mux_v
    port map (
            O => \N__29041\,
            I => \N__29000\
        );

    \I__6368\ : Span4Mux_h
    port map (
            O => \N__29036\,
            I => \N__29000\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__29027\,
            I => \N__29000\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__29024\,
            I => cmd_12
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__29021\,
            I => cmd_12
        );

    \I__6364\ : Odrv12
    port map (
            O => \N__29018\,
            I => cmd_12
        );

    \I__6363\ : Odrv4
    port map (
            O => \N__29015\,
            I => cmd_12
        );

    \I__6362\ : Odrv4
    port map (
            O => \N__29012\,
            I => cmd_12
        );

    \I__6361\ : Odrv4
    port map (
            O => \N__29007\,
            I => cmd_12
        );

    \I__6360\ : Odrv4
    port map (
            O => \N__29000\,
            I => cmd_12
        );

    \I__6359\ : CascadeMux
    port map (
            O => \N__28985\,
            I => \N__28982\
        );

    \I__6358\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28979\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__28979\,
            I => \N__28975\
        );

    \I__6356\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28972\
        );

    \I__6355\ : Span4Mux_h
    port map (
            O => \N__28975\,
            I => \N__28969\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__28972\,
            I => fwd_7
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__28969\,
            I => fwd_7
        );

    \I__6352\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28958\
        );

    \I__6351\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28958\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__28958\,
            I => \N__28951\
        );

    \I__6349\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28946\
        );

    \I__6348\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28946\
        );

    \I__6347\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28941\
        );

    \I__6346\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28941\
        );

    \I__6345\ : Span4Mux_v
    port map (
            O => \N__28951\,
            I => \N__28938\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__28946\,
            I => \N__28935\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__28941\,
            I => \Inst_core.Inst_trigger.levelReg_0\
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__28938\,
            I => \Inst_core.Inst_trigger.levelReg_0\
        );

    \I__6341\ : Odrv4
    port map (
            O => \N__28935\,
            I => \Inst_core.Inst_trigger.levelReg_0\
        );

    \I__6340\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28924\
        );

    \I__6339\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28921\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__28924\,
            I => \N__28918\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__28921\,
            I => \configRegister_17_adj_1343\
        );

    \I__6336\ : Odrv4
    port map (
            O => \N__28918\,
            I => \configRegister_17_adj_1343\
        );

    \I__6335\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28904\
        );

    \I__6334\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28904\
        );

    \I__6333\ : InMux
    port map (
            O => \N__28911\,
            I => \N__28899\
        );

    \I__6332\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28899\
        );

    \I__6331\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28896\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__28904\,
            I => \N__28893\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__28899\,
            I => \N__28890\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__28896\,
            I => \N__28885\
        );

    \I__6327\ : Span4Mux_v
    port map (
            O => \N__28893\,
            I => \N__28885\
        );

    \I__6326\ : Odrv4
    port map (
            O => \N__28890\,
            I => \Inst_core.Inst_trigger.levelReg_1\
        );

    \I__6325\ : Odrv4
    port map (
            O => \N__28885\,
            I => \Inst_core.Inst_trigger.levelReg_1\
        );

    \I__6324\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28874\
        );

    \I__6323\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28874\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28871\
        );

    \I__6321\ : Span12Mux_s5_v
    port map (
            O => \N__28871\,
            I => \N__28868\
        );

    \I__6320\ : Odrv12
    port map (
            O => \N__28868\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n99\
        );

    \I__6319\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28862\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__28862\,
            I => \N__28858\
        );

    \I__6317\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28855\
        );

    \I__6316\ : Odrv12
    port map (
            O => \N__28858\,
            I => \valueRegister_4_adj_1372\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__28855\,
            I => \valueRegister_4_adj_1372\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__28850\,
            I => \N__28847\
        );

    \I__6313\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28840\
        );

    \I__6311\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28837\
        );

    \I__6310\ : Odrv12
    port map (
            O => \N__28840\,
            I => \configRegister_15_adj_1305\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__28837\,
            I => \configRegister_15_adj_1305\
        );

    \I__6308\ : CascadeMux
    port map (
            O => \N__28832\,
            I => \N__28829\
        );

    \I__6307\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28826\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__28826\,
            I => \N__28822\
        );

    \I__6305\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28819\
        );

    \I__6304\ : Span4Mux_h
    port map (
            O => \N__28822\,
            I => \N__28816\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__28819\,
            I => bwd_15
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__28816\,
            I => bwd_15
        );

    \I__6301\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28808\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__28808\,
            I => \N__28805\
        );

    \I__6299\ : Span4Mux_v
    port map (
            O => \N__28805\,
            I => \N__28801\
        );

    \I__6298\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28798\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__28801\,
            I => \configRegister_13_adj_1307\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__28798\,
            I => \configRegister_13_adj_1307\
        );

    \I__6295\ : InMux
    port map (
            O => \N__28793\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7896\
        );

    \I__6294\ : CascadeMux
    port map (
            O => \N__28790\,
            I => \N__28786\
        );

    \I__6293\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28783\
        );

    \I__6292\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28780\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__28783\,
            I => \N__28777\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__28780\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__28777\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14\
        );

    \I__6288\ : InMux
    port map (
            O => \N__28772\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7897\
        );

    \I__6287\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28763\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__28768\,
            I => \N__28758\
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__28767\,
            I => \N__28754\
        );

    \I__6284\ : CascadeMux
    port map (
            O => \N__28766\,
            I => \N__28750\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__28763\,
            I => \N__28746\
        );

    \I__6282\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28726\
        );

    \I__6281\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28726\
        );

    \I__6280\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28726\
        );

    \I__6279\ : InMux
    port map (
            O => \N__28757\,
            I => \N__28726\
        );

    \I__6278\ : InMux
    port map (
            O => \N__28754\,
            I => \N__28726\
        );

    \I__6277\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28726\
        );

    \I__6276\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28726\
        );

    \I__6275\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28726\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__28746\,
            I => \N__28723\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__28745\,
            I => \N__28719\
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__28744\,
            I => \N__28715\
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__28743\,
            I => \N__28711\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__28726\,
            I => \N__28705\
        );

    \I__6269\ : Span4Mux_v
    port map (
            O => \N__28723\,
            I => \N__28705\
        );

    \I__6268\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28690\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28690\
        );

    \I__6266\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28690\
        );

    \I__6265\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28690\
        );

    \I__6264\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28690\
        );

    \I__6263\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28690\
        );

    \I__6262\ : InMux
    port map (
            O => \N__28710\,
            I => \N__28690\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__28705\,
            I => \N__28687\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__28690\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n1662\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__28687\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n1662\
        );

    \I__6258\ : InMux
    port map (
            O => \N__28682\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7898\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__28679\,
            I => \N__28676\
        );

    \I__6256\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28672\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28669\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__28672\,
            I => \N__28666\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__28669\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__28666\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15\
        );

    \I__6251\ : CEMux
    port map (
            O => \N__28661\,
            I => \N__28658\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28654\
        );

    \I__6249\ : CEMux
    port map (
            O => \N__28657\,
            I => \N__28651\
        );

    \I__6248\ : Odrv12
    port map (
            O => \N__28654\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4144\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__28651\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4144\
        );

    \I__6246\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28643\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__28643\,
            I => \N__28639\
        );

    \I__6244\ : CascadeMux
    port map (
            O => \N__28642\,
            I => \N__28636\
        );

    \I__6243\ : Span4Mux_v
    port map (
            O => \N__28639\,
            I => \N__28632\
        );

    \I__6242\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28627\
        );

    \I__6241\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28627\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__28632\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__28627\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2\
        );

    \I__6238\ : SRMux
    port map (
            O => \N__28622\,
            I => \N__28619\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__28619\,
            I => \N__28616\
        );

    \I__6236\ : Span4Mux_s2_h
    port map (
            O => \N__28616\,
            I => \N__28613\
        );

    \I__6235\ : Span4Mux_h
    port map (
            O => \N__28613\,
            I => \N__28610\
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__28610\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4761\
        );

    \I__6233\ : CascadeMux
    port map (
            O => \N__28607\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n2_cascade_\
        );

    \I__6232\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28601\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28598\
        );

    \I__6230\ : Span4Mux_v
    port map (
            O => \N__28598\,
            I => \N__28595\
        );

    \I__6229\ : Sp12to4
    port map (
            O => \N__28595\,
            I => \N__28592\
        );

    \I__6228\ : Odrv12
    port map (
            O => \N__28592\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register\
        );

    \I__6227\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__28586\,
            I => \N__28583\
        );

    \I__6225\ : Span4Mux_v
    port map (
            O => \N__28583\,
            I => \N__28580\
        );

    \I__6224\ : Odrv4
    port map (
            O => \N__28580\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n100\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__28577\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n100_cascade_\
        );

    \I__6222\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28570\
        );

    \I__6221\ : CascadeMux
    port map (
            O => \N__28573\,
            I => \N__28567\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__28570\,
            I => \N__28564\
        );

    \I__6219\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28561\
        );

    \I__6218\ : Span4Mux_s2_h
    port map (
            O => \N__28564\,
            I => \N__28558\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__28561\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n450\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__28558\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n450\
        );

    \I__6215\ : InMux
    port map (
            O => \N__28553\,
            I => \N__28550\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__28550\,
            I => \N__28546\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28543\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__28546\,
            I => \configRegister_5_adj_1315\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__28543\,
            I => \configRegister_5_adj_1315\
        );

    \I__6210\ : InMux
    port map (
            O => \N__28538\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7888\
        );

    \I__6209\ : InMux
    port map (
            O => \N__28535\,
            I => \N__28532\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__28532\,
            I => \N__28528\
        );

    \I__6207\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28525\
        );

    \I__6206\ : Odrv4
    port map (
            O => \N__28528\,
            I => \configRegister_6_adj_1314\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__28525\,
            I => \configRegister_6_adj_1314\
        );

    \I__6204\ : InMux
    port map (
            O => \N__28520\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7889\
        );

    \I__6203\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__6201\ : Span4Mux_v
    port map (
            O => \N__28511\,
            I => \N__28508\
        );

    \I__6200\ : Span4Mux_s1_h
    port map (
            O => \N__28508\,
            I => \N__28504\
        );

    \I__6199\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28501\
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__28504\,
            I => \configRegister_7_adj_1313\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__28501\,
            I => \configRegister_7_adj_1313\
        );

    \I__6196\ : InMux
    port map (
            O => \N__28496\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7890\
        );

    \I__6195\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28490\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28486\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__28489\,
            I => \N__28483\
        );

    \I__6192\ : Span12Mux_s5_h
    port map (
            O => \N__28486\,
            I => \N__28480\
        );

    \I__6191\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28477\
        );

    \I__6190\ : Odrv12
    port map (
            O => \N__28480\,
            I => \configRegister_8_adj_1312\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__28477\,
            I => \configRegister_8_adj_1312\
        );

    \I__6188\ : InMux
    port map (
            O => \N__28472\,
            I => \bfn_11_5_0_\
        );

    \I__6187\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__28466\,
            I => \N__28463\
        );

    \I__6185\ : Span4Mux_s2_h
    port map (
            O => \N__28463\,
            I => \N__28459\
        );

    \I__6184\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28456\
        );

    \I__6183\ : Odrv4
    port map (
            O => \N__28459\,
            I => \configRegister_9_adj_1311\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__28456\,
            I => \configRegister_9_adj_1311\
        );

    \I__6181\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28447\
        );

    \I__6180\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28444\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__28447\,
            I => \N__28441\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__28444\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9\
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__28441\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9\
        );

    \I__6176\ : InMux
    port map (
            O => \N__28436\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7892\
        );

    \I__6175\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28427\
        );

    \I__6173\ : Span4Mux_v
    port map (
            O => \N__28427\,
            I => \N__28423\
        );

    \I__6172\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28420\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__28423\,
            I => \configRegister_10_adj_1310\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__28420\,
            I => \configRegister_10_adj_1310\
        );

    \I__6169\ : InMux
    port map (
            O => \N__28415\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7893\
        );

    \I__6168\ : InMux
    port map (
            O => \N__28412\,
            I => \N__28409\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__28409\,
            I => \N__28406\
        );

    \I__6166\ : Span4Mux_h
    port map (
            O => \N__28406\,
            I => \N__28402\
        );

    \I__6165\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28399\
        );

    \I__6164\ : Odrv4
    port map (
            O => \N__28402\,
            I => \configRegister_11_adj_1309\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__28399\,
            I => \configRegister_11_adj_1309\
        );

    \I__6162\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28390\
        );

    \I__6161\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28387\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__28390\,
            I => \N__28384\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__28387\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__28384\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11\
        );

    \I__6157\ : InMux
    port map (
            O => \N__28379\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7894\
        );

    \I__6156\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28373\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__28373\,
            I => \N__28369\
        );

    \I__6154\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28366\
        );

    \I__6153\ : Odrv12
    port map (
            O => \N__28369\,
            I => \configRegister_12_adj_1308\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__28366\,
            I => \configRegister_12_adj_1308\
        );

    \I__6151\ : InMux
    port map (
            O => \N__28361\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7895\
        );

    \I__6150\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__28355\,
            I => \N__28352\
        );

    \I__6148\ : Span4Mux_s2_v
    port map (
            O => \N__28352\,
            I => \N__28348\
        );

    \I__6147\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__28348\,
            I => \Inst_core.n8837\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__28345\,
            I => \Inst_core.n8837\
        );

    \I__6144\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__6143\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28327\
        );

    \I__6142\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28327\
        );

    \I__6141\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28327\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28321\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__28327\,
            I => \N__28321\
        );

    \I__6138\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28318\
        );

    \I__6137\ : Span4Mux_v
    port map (
            O => \N__28321\,
            I => \N__28315\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__28318\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.state_1\
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__28315\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.state_1\
        );

    \I__6134\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28306\
        );

    \I__6133\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28303\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__28306\,
            I => \N__28300\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__28303\,
            I => \configRegister_0_adj_1320\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__28300\,
            I => \configRegister_0_adj_1320\
        );

    \I__6129\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__28292\,
            I => \N__28289\
        );

    \I__6127\ : Span4Mux_s2_h
    port map (
            O => \N__28289\,
            I => \N__28286\
        );

    \I__6126\ : Span4Mux_v
    port map (
            O => \N__28286\,
            I => \N__28283\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__28283\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9055\
        );

    \I__6124\ : InMux
    port map (
            O => \N__28280\,
            I => \bfn_11_4_0_\
        );

    \I__6123\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28274\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__28274\,
            I => \N__28271\
        );

    \I__6121\ : Span4Mux_s1_h
    port map (
            O => \N__28271\,
            I => \N__28267\
        );

    \I__6120\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28264\
        );

    \I__6119\ : Odrv4
    port map (
            O => \N__28267\,
            I => \configRegister_1_adj_1319\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__28264\,
            I => \configRegister_1_adj_1319\
        );

    \I__6117\ : InMux
    port map (
            O => \N__28259\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7884\
        );

    \I__6116\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28252\
        );

    \I__6115\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28249\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__28252\,
            I => \N__28246\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__28249\,
            I => \configRegister_2_adj_1318\
        );

    \I__6112\ : Odrv4
    port map (
            O => \N__28246\,
            I => \configRegister_2_adj_1318\
        );

    \I__6111\ : InMux
    port map (
            O => \N__28241\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7885\
        );

    \I__6110\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28235\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__28235\,
            I => \N__28231\
        );

    \I__6108\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28228\
        );

    \I__6107\ : Odrv4
    port map (
            O => \N__28231\,
            I => \configRegister_3_adj_1317\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__28228\,
            I => \configRegister_3_adj_1317\
        );

    \I__6105\ : InMux
    port map (
            O => \N__28223\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7886\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28217\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__28217\,
            I => \N__28214\
        );

    \I__6102\ : Span4Mux_s3_h
    port map (
            O => \N__28214\,
            I => \N__28210\
        );

    \I__6101\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28207\
        );

    \I__6100\ : Odrv4
    port map (
            O => \N__28210\,
            I => \configRegister_4_adj_1316\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__28207\,
            I => \configRegister_4_adj_1316\
        );

    \I__6098\ : InMux
    port map (
            O => \N__28202\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7887\
        );

    \I__6097\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28196\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__28196\,
            I => \N__28193\
        );

    \I__6095\ : Span4Mux_s3_v
    port map (
            O => \N__28193\,
            I => \N__28187\
        );

    \I__6094\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28184\
        );

    \I__6093\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28179\
        );

    \I__6092\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28179\
        );

    \I__6091\ : Span4Mux_h
    port map (
            O => \N__28187\,
            I => \N__28171\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__28184\,
            I => \N__28171\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__28179\,
            I => \N__28168\
        );

    \I__6088\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28165\
        );

    \I__6087\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28162\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__28176\,
            I => \N__28159\
        );

    \I__6085\ : Span4Mux_v
    port map (
            O => \N__28171\,
            I => \N__28156\
        );

    \I__6084\ : Span12Mux_s4_h
    port map (
            O => \N__28168\,
            I => \N__28151\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__28165\,
            I => \N__28151\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__28162\,
            I => \N__28148\
        );

    \I__6081\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28145\
        );

    \I__6080\ : Odrv4
    port map (
            O => \N__28156\,
            I => cmd_35
        );

    \I__6079\ : Odrv12
    port map (
            O => \N__28151\,
            I => cmd_35
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__28148\,
            I => cmd_35
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__28145\,
            I => cmd_35
        );

    \I__6076\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28133\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28129\
        );

    \I__6074\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__28129\,
            I => \configRegister_0_adj_1360\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__28126\,
            I => \configRegister_0_adj_1360\
        );

    \I__6071\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28117\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__28120\,
            I => \N__28114\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__28117\,
            I => \N__28110\
        );

    \I__6068\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28105\
        );

    \I__6067\ : InMux
    port map (
            O => \N__28113\,
            I => \N__28105\
        );

    \I__6066\ : Span4Mux_h
    port map (
            O => \N__28110\,
            I => \N__28102\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__28105\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__28102\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__6062\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__28091\,
            I => \N__28088\
        );

    \I__6060\ : Span4Mux_s3_h
    port map (
            O => \N__28088\,
            I => \N__28082\
        );

    \I__6059\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28078\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__28086\,
            I => \N__28073\
        );

    \I__6057\ : InMux
    port map (
            O => \N__28085\,
            I => \N__28069\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__28082\,
            I => \N__28066\
        );

    \I__6055\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28063\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__28078\,
            I => \N__28060\
        );

    \I__6053\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28057\
        );

    \I__6052\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28054\
        );

    \I__6051\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28051\
        );

    \I__6050\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28048\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28045\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__28066\,
            I => \N__28040\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__28063\,
            I => \N__28040\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__28060\,
            I => \N__28037\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28034\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__28054\,
            I => \N__28029\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__28051\,
            I => \N__28029\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__28048\,
            I => \N__28024\
        );

    \I__6041\ : Span4Mux_h
    port map (
            O => \N__28045\,
            I => \N__28019\
        );

    \I__6040\ : Span4Mux_v
    port map (
            O => \N__28040\,
            I => \N__28019\
        );

    \I__6039\ : Span4Mux_h
    port map (
            O => \N__28037\,
            I => \N__28012\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__28034\,
            I => \N__28012\
        );

    \I__6037\ : Span4Mux_h
    port map (
            O => \N__28029\,
            I => \N__28012\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28009\
        );

    \I__6035\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28006\
        );

    \I__6034\ : Span4Mux_v
    port map (
            O => \N__28024\,
            I => \N__28001\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__28019\,
            I => \N__28001\
        );

    \I__6032\ : Span4Mux_v
    port map (
            O => \N__28012\,
            I => \N__27998\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__28009\,
            I => \N__27995\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__28006\,
            I => \memoryOut_4\
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__28001\,
            I => \memoryOut_4\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__27998\,
            I => \memoryOut_4\
        );

    \I__6027\ : Odrv12
    port map (
            O => \N__27995\,
            I => \memoryOut_4\
        );

    \I__6026\ : SRMux
    port map (
            O => \N__27986\,
            I => \N__27983\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__27983\,
            I => \N__27980\
        );

    \I__6024\ : Span4Mux_s3_v
    port map (
            O => \N__27980\,
            I => \N__27977\
        );

    \I__6023\ : Span4Mux_s1_h
    port map (
            O => \N__27977\,
            I => \N__27974\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__27974\,
            I => \N__27971\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__27971\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4763\
        );

    \I__6020\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__6018\ : Span4Mux_s2_h
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__27959\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_5\
        );

    \I__6016\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__27953\,
            I => \N__27950\
        );

    \I__6014\ : Odrv12
    port map (
            O => \N__27950\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_7\
        );

    \I__6013\ : CascadeMux
    port map (
            O => \N__27947\,
            I => \N__27944\
        );

    \I__6012\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27941\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__27941\,
            I => \N__27938\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__27938\,
            I => \N__27935\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__27935\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_6\
        );

    \I__6008\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27929\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__27929\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_4\
        );

    \I__6006\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27923\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27920\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__27920\,
            I => \N__27917\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__27917\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n11\
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__27914\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n6675_cascade_\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__27911\,
            I => \N__27907\
        );

    \I__6000\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27904\
        );

    \I__5999\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27901\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__27904\,
            I => \N__27898\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27901\,
            I => \N__27895\
        );

    \I__5996\ : Span4Mux_v
    port map (
            O => \N__27898\,
            I => \N__27892\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__27895\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n564\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__27892\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n564\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__27887\,
            I => \N__27884\
        );

    \I__5992\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27881\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__27881\,
            I => \N__27877\
        );

    \I__5990\ : InMux
    port map (
            O => \N__27880\,
            I => \N__27873\
        );

    \I__5989\ : Span4Mux_v
    port map (
            O => \N__27877\,
            I => \N__27870\
        );

    \I__5988\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27867\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__27873\,
            I => \Inst_core.Inst_sampler.counter_17\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__27870\,
            I => \Inst_core.Inst_sampler.counter_17\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__27867\,
            I => \Inst_core.Inst_sampler.counter_17\
        );

    \I__5984\ : InMux
    port map (
            O => \N__27860\,
            I => \Inst_core.Inst_sampler.n7964\
        );

    \I__5983\ : InMux
    port map (
            O => \N__27857\,
            I => \Inst_core.Inst_sampler.n7965\
        );

    \I__5982\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27851\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__27851\,
            I => \N__27846\
        );

    \I__5980\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27843\
        );

    \I__5979\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27840\
        );

    \I__5978\ : Span4Mux_h
    port map (
            O => \N__27846\,
            I => \N__27837\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__27843\,
            I => \N__27834\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__27840\,
            I => \Inst_core.Inst_sampler.counter_19\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__27837\,
            I => \Inst_core.Inst_sampler.counter_19\
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__27834\,
            I => \Inst_core.Inst_sampler.counter_19\
        );

    \I__5973\ : InMux
    port map (
            O => \N__27827\,
            I => \Inst_core.Inst_sampler.n7966\
        );

    \I__5972\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27819\
        );

    \I__5971\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27814\
        );

    \I__5970\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27814\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__27819\,
            I => \Inst_core.Inst_sampler.counter_20\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__27814\,
            I => \Inst_core.Inst_sampler.counter_20\
        );

    \I__5967\ : InMux
    port map (
            O => \N__27809\,
            I => \Inst_core.Inst_sampler.n7967\
        );

    \I__5966\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27802\
        );

    \I__5965\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27799\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__27802\,
            I => \N__27795\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27792\
        );

    \I__5962\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27789\
        );

    \I__5961\ : Span4Mux_v
    port map (
            O => \N__27795\,
            I => \N__27786\
        );

    \I__5960\ : Span4Mux_v
    port map (
            O => \N__27792\,
            I => \N__27783\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__27789\,
            I => \Inst_core.Inst_sampler.counter_21\
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__27786\,
            I => \Inst_core.Inst_sampler.counter_21\
        );

    \I__5957\ : Odrv4
    port map (
            O => \N__27783\,
            I => \Inst_core.Inst_sampler.counter_21\
        );

    \I__5956\ : InMux
    port map (
            O => \N__27776\,
            I => \Inst_core.Inst_sampler.n7968\
        );

    \I__5955\ : InMux
    port map (
            O => \N__27773\,
            I => \Inst_core.Inst_sampler.n7969\
        );

    \I__5954\ : InMux
    port map (
            O => \N__27770\,
            I => \Inst_core.Inst_sampler.n7970\
        );

    \I__5953\ : SRMux
    port map (
            O => \N__27767\,
            I => \N__27764\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__27764\,
            I => \N__27760\
        );

    \I__5951\ : SRMux
    port map (
            O => \N__27763\,
            I => \N__27757\
        );

    \I__5950\ : Span4Mux_s1_v
    port map (
            O => \N__27760\,
            I => \N__27751\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__27757\,
            I => \N__27751\
        );

    \I__5948\ : SRMux
    port map (
            O => \N__27756\,
            I => \N__27748\
        );

    \I__5947\ : Span4Mux_v
    port map (
            O => \N__27751\,
            I => \N__27745\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__27748\,
            I => \N__27742\
        );

    \I__5945\ : Span4Mux_s3_h
    port map (
            O => \N__27745\,
            I => \N__27737\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__27742\,
            I => \N__27737\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__27737\,
            I => \N__27734\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__27734\,
            I => \N__27731\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__27731\,
            I => \Inst_core.Inst_sampler.n1700\
        );

    \I__5940\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27725\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__27725\,
            I => \N__27720\
        );

    \I__5938\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27715\
        );

    \I__5937\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27715\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__27720\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__27715\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997\
        );

    \I__5934\ : SRMux
    port map (
            O => \N__27710\,
            I => \N__27707\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__5932\ : Odrv12
    port map (
            O => \N__27704\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n8622\
        );

    \I__5931\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27696\
        );

    \I__5930\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27693\
        );

    \I__5929\ : InMux
    port map (
            O => \N__27699\,
            I => \N__27690\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__27696\,
            I => \N__27687\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__27693\,
            I => \Inst_core.Inst_sampler.counter_9\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__27690\,
            I => \Inst_core.Inst_sampler.counter_9\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__27687\,
            I => \Inst_core.Inst_sampler.counter_9\
        );

    \I__5924\ : InMux
    port map (
            O => \N__27680\,
            I => \Inst_core.Inst_sampler.n7956\
        );

    \I__5923\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27670\
        );

    \I__5922\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27670\
        );

    \I__5921\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27667\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__27670\,
            I => \N__27664\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__27667\,
            I => \Inst_core.Inst_sampler.counter_10\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__27664\,
            I => \Inst_core.Inst_sampler.counter_10\
        );

    \I__5917\ : InMux
    port map (
            O => \N__27659\,
            I => \Inst_core.Inst_sampler.n7957\
        );

    \I__5916\ : InMux
    port map (
            O => \N__27656\,
            I => \Inst_core.Inst_sampler.n7958\
        );

    \I__5915\ : InMux
    port map (
            O => \N__27653\,
            I => \Inst_core.Inst_sampler.n7959\
        );

    \I__5914\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27645\
        );

    \I__5913\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27640\
        );

    \I__5912\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27640\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__27645\,
            I => \Inst_core.Inst_sampler.counter_13\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__27640\,
            I => \Inst_core.Inst_sampler.counter_13\
        );

    \I__5909\ : InMux
    port map (
            O => \N__27635\,
            I => \Inst_core.Inst_sampler.n7960\
        );

    \I__5908\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27627\
        );

    \I__5907\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27622\
        );

    \I__5906\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27622\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__27627\,
            I => \Inst_core.Inst_sampler.counter_14\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__27622\,
            I => \Inst_core.Inst_sampler.counter_14\
        );

    \I__5903\ : InMux
    port map (
            O => \N__27617\,
            I => \Inst_core.Inst_sampler.n7961\
        );

    \I__5902\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27609\
        );

    \I__5901\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27604\
        );

    \I__5900\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27604\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__27609\,
            I => \Inst_core.Inst_sampler.counter_15\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__27604\,
            I => \Inst_core.Inst_sampler.counter_15\
        );

    \I__5897\ : InMux
    port map (
            O => \N__27599\,
            I => \Inst_core.Inst_sampler.n7962\
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__27596\,
            I => \N__27593\
        );

    \I__5895\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27588\
        );

    \I__5894\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27585\
        );

    \I__5893\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27582\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27579\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__27585\,
            I => \N__27576\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__27582\,
            I => \Inst_core.Inst_sampler.counter_16\
        );

    \I__5889\ : Odrv12
    port map (
            O => \N__27579\,
            I => \Inst_core.Inst_sampler.counter_16\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__27576\,
            I => \Inst_core.Inst_sampler.counter_16\
        );

    \I__5887\ : InMux
    port map (
            O => \N__27569\,
            I => \bfn_9_16_0_\
        );

    \I__5886\ : InMux
    port map (
            O => \N__27566\,
            I => \bfn_9_14_0_\
        );

    \I__5885\ : InMux
    port map (
            O => \N__27563\,
            I => \Inst_core.Inst_sampler.n7948\
        );

    \I__5884\ : InMux
    port map (
            O => \N__27560\,
            I => \Inst_core.Inst_sampler.n7949\
        );

    \I__5883\ : InMux
    port map (
            O => \N__27557\,
            I => \Inst_core.Inst_sampler.n7950\
        );

    \I__5882\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27549\
        );

    \I__5881\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27546\
        );

    \I__5880\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27543\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__27549\,
            I => \Inst_core.Inst_sampler.counter_4\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__27546\,
            I => \Inst_core.Inst_sampler.counter_4\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__27543\,
            I => \Inst_core.Inst_sampler.counter_4\
        );

    \I__5876\ : InMux
    port map (
            O => \N__27536\,
            I => \Inst_core.Inst_sampler.n7951\
        );

    \I__5875\ : InMux
    port map (
            O => \N__27533\,
            I => \Inst_core.Inst_sampler.n7952\
        );

    \I__5874\ : InMux
    port map (
            O => \N__27530\,
            I => \Inst_core.Inst_sampler.n7953\
        );

    \I__5873\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27522\
        );

    \I__5872\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27519\
        );

    \I__5871\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27516\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__27522\,
            I => \Inst_core.Inst_sampler.counter_7\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__27519\,
            I => \Inst_core.Inst_sampler.counter_7\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__27516\,
            I => \Inst_core.Inst_sampler.counter_7\
        );

    \I__5867\ : InMux
    port map (
            O => \N__27509\,
            I => \Inst_core.Inst_sampler.n7954\
        );

    \I__5866\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27503\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__27503\,
            I => \N__27498\
        );

    \I__5864\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27495\
        );

    \I__5863\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27492\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__27498\,
            I => \N__27489\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27486\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__27492\,
            I => \Inst_core.Inst_sampler.counter_8\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__27489\,
            I => \Inst_core.Inst_sampler.counter_8\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__27486\,
            I => \Inst_core.Inst_sampler.counter_8\
        );

    \I__5857\ : InMux
    port map (
            O => \N__27479\,
            I => \bfn_9_15_0_\
        );

    \I__5856\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27472\
        );

    \I__5855\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27469\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__27472\,
            I => \maskRegister_1_adj_1327\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__27469\,
            I => \maskRegister_1_adj_1327\
        );

    \I__5852\ : SRMux
    port map (
            O => \N__27464\,
            I => \N__27461\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__27461\,
            I => \N__27458\
        );

    \I__5850\ : Span4Mux_v
    port map (
            O => \N__27458\,
            I => \N__27455\
        );

    \I__5849\ : Sp12to4
    port map (
            O => \N__27455\,
            I => \N__27452\
        );

    \I__5848\ : Odrv12
    port map (
            O => \N__27452\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4753\
        );

    \I__5847\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27445\
        );

    \I__5846\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27442\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__27445\,
            I => \maskRegister_2_adj_1326\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__27442\,
            I => \maskRegister_2_adj_1326\
        );

    \I__5843\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27433\
        );

    \I__5842\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27430\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__27433\,
            I => \N__27427\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__27430\,
            I => \maskRegister_3_adj_1325\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__27427\,
            I => \maskRegister_3_adj_1325\
        );

    \I__5838\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27419\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__27419\,
            I => \N__27416\
        );

    \I__5836\ : Span4Mux_s3_h
    port map (
            O => \N__27416\,
            I => \N__27412\
        );

    \I__5835\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27409\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__27412\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__27409\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6\
        );

    \I__5832\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__27401\,
            I => \N__27398\
        );

    \I__5830\ : Span4Mux_v
    port map (
            O => \N__27398\,
            I => \N__27395\
        );

    \I__5829\ : Span4Mux_v
    port map (
            O => \N__27395\,
            I => \N__27391\
        );

    \I__5828\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27388\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__27391\,
            I => \valueRegister_6_adj_1330\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__27388\,
            I => \valueRegister_6_adj_1330\
        );

    \I__5825\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27380\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__27380\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_6\
        );

    \I__5823\ : SRMux
    port map (
            O => \N__27377\,
            I => \N__27374\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__27374\,
            I => \N__27371\
        );

    \I__5821\ : Span4Mux_v
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__5820\ : Span4Mux_s2_h
    port map (
            O => \N__27368\,
            I => \N__27365\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__27365\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4758\
        );

    \I__5818\ : InMux
    port map (
            O => \N__27362\,
            I => \N__27357\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__27361\,
            I => \N__27354\
        );

    \I__5816\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27351\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__27357\,
            I => \N__27348\
        );

    \I__5814\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27345\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__27351\,
            I => \N__27340\
        );

    \I__5812\ : Span4Mux_h
    port map (
            O => \N__27348\,
            I => \N__27340\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27337\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__27340\,
            I => divider_4
        );

    \I__5809\ : Odrv12
    port map (
            O => \N__27337\,
            I => divider_4
        );

    \I__5808\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__27329\,
            I => \Inst_core.Inst_sampler.n30\
        );

    \I__5806\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27323\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27320\
        );

    \I__5804\ : Odrv4
    port map (
            O => \N__27320\,
            I => \Inst_core.Inst_sampler.n8592\
        );

    \I__5803\ : InMux
    port map (
            O => \N__27317\,
            I => \N__27310\
        );

    \I__5802\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27310\
        );

    \I__5801\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27307\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__27310\,
            I => \N__27304\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__27307\,
            I => divider_2
        );

    \I__5798\ : Odrv12
    port map (
            O => \N__27304\,
            I => divider_2
        );

    \I__5797\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27291\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27288\
        );

    \I__5794\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27285\
        );

    \I__5793\ : Sp12to4
    port map (
            O => \N__27291\,
            I => \N__27280\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__27288\,
            I => \N__27280\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__27285\,
            I => divider_10
        );

    \I__5790\ : Odrv12
    port map (
            O => \N__27280\,
            I => divider_10
        );

    \I__5789\ : CascadeMux
    port map (
            O => \N__27275\,
            I => \N__27271\
        );

    \I__5788\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27266\
        );

    \I__5787\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27266\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27263\
        );

    \I__5785\ : Span4Mux_h
    port map (
            O => \N__27263\,
            I => \N__27259\
        );

    \I__5784\ : InMux
    port map (
            O => \N__27262\,
            I => \N__27256\
        );

    \I__5783\ : Span4Mux_v
    port map (
            O => \N__27259\,
            I => \N__27253\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__27256\,
            I => divider_8
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__27253\,
            I => divider_8
        );

    \I__5780\ : CascadeMux
    port map (
            O => \N__27248\,
            I => \N__27244\
        );

    \I__5779\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27241\
        );

    \I__5778\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27238\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__27241\,
            I => \N__27234\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__27238\,
            I => \N__27231\
        );

    \I__5775\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27228\
        );

    \I__5774\ : Span4Mux_v
    port map (
            O => \N__27234\,
            I => \N__27225\
        );

    \I__5773\ : Span12Mux_s6_v
    port map (
            O => \N__27231\,
            I => \N__27222\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__27228\,
            I => divider_17
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__27225\,
            I => divider_17
        );

    \I__5770\ : Odrv12
    port map (
            O => \N__27222\,
            I => divider_17
        );

    \I__5769\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__27212\,
            I => \Inst_core.Inst_sampler.n8588\
        );

    \I__5767\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27202\
        );

    \I__5766\ : CascadeMux
    port map (
            O => \N__27208\,
            I => \N__27194\
        );

    \I__5765\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27188\
        );

    \I__5764\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27183\
        );

    \I__5763\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27183\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__27202\,
            I => \N__27180\
        );

    \I__5761\ : InMux
    port map (
            O => \N__27201\,
            I => \N__27175\
        );

    \I__5760\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27175\
        );

    \I__5759\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27171\
        );

    \I__5758\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27168\
        );

    \I__5757\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27165\
        );

    \I__5756\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27162\
        );

    \I__5755\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27159\
        );

    \I__5754\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27156\
        );

    \I__5753\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27153\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__27188\,
            I => \N__27150\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__27183\,
            I => \N__27143\
        );

    \I__5750\ : Span4Mux_s3_v
    port map (
            O => \N__27180\,
            I => \N__27143\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__27175\,
            I => \N__27143\
        );

    \I__5748\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27137\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27134\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__27168\,
            I => \N__27129\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__27165\,
            I => \N__27129\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__27162\,
            I => \N__27124\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__27159\,
            I => \N__27124\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__27156\,
            I => \N__27121\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__27153\,
            I => \N__27114\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__27150\,
            I => \N__27114\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__27143\,
            I => \N__27114\
        );

    \I__5738\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27107\
        );

    \I__5737\ : InMux
    port map (
            O => \N__27141\,
            I => \N__27107\
        );

    \I__5736\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27107\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__27137\,
            I => \N__27104\
        );

    \I__5734\ : Span4Mux_v
    port map (
            O => \N__27134\,
            I => \N__27101\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__27129\,
            I => \N__27098\
        );

    \I__5732\ : Span4Mux_h
    port map (
            O => \N__27124\,
            I => \N__27095\
        );

    \I__5731\ : Span4Mux_h
    port map (
            O => \N__27121\,
            I => \N__27090\
        );

    \I__5730\ : Span4Mux_h
    port map (
            O => \N__27114\,
            I => \N__27090\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__27107\,
            I => cmd_15
        );

    \I__5728\ : Odrv4
    port map (
            O => \N__27104\,
            I => cmd_15
        );

    \I__5727\ : Odrv4
    port map (
            O => \N__27101\,
            I => cmd_15
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__27098\,
            I => cmd_15
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__27095\,
            I => cmd_15
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__27090\,
            I => cmd_15
        );

    \I__5723\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27073\
        );

    \I__5722\ : InMux
    port map (
            O => \N__27076\,
            I => \N__27070\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__27073\,
            I => bwd_7
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__27070\,
            I => bwd_7
        );

    \I__5719\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27061\
        );

    \I__5718\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27058\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__27061\,
            I => fwd_10
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__27058\,
            I => fwd_10
        );

    \I__5715\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27044\
        );

    \I__5714\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27044\
        );

    \I__5713\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27039\
        );

    \I__5712\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27036\
        );

    \I__5711\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27033\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__27044\,
            I => \N__27030\
        );

    \I__5709\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27027\
        );

    \I__5708\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27024\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__27018\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__27036\,
            I => \N__27018\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__27033\,
            I => \N__27015\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__27030\,
            I => \N__27008\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__27008\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27008\
        );

    \I__5701\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27005\
        );

    \I__5700\ : Span4Mux_h
    port map (
            O => \N__27018\,
            I => \N__27002\
        );

    \I__5699\ : Span4Mux_s3_h
    port map (
            O => \N__27015\,
            I => \N__26997\
        );

    \I__5698\ : Span4Mux_v
    port map (
            O => \N__27008\,
            I => \N__26997\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__27005\,
            I => \N__26994\
        );

    \I__5696\ : Span4Mux_v
    port map (
            O => \N__27002\,
            I => \N__26991\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__26997\,
            I => \N__26988\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__26994\,
            I => wrtrigmask_2
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__26991\,
            I => wrtrigmask_2
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__26988\,
            I => wrtrigmask_2
        );

    \I__5691\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26977\
        );

    \I__5690\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26974\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__26977\,
            I => \maskRegister_4_adj_1324\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__26974\,
            I => \maskRegister_4_adj_1324\
        );

    \I__5687\ : CascadeMux
    port map (
            O => \N__26969\,
            I => \N__26966\
        );

    \I__5686\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26963\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__26963\,
            I => \N__26959\
        );

    \I__5684\ : InMux
    port map (
            O => \N__26962\,
            I => \N__26956\
        );

    \I__5683\ : Span4Mux_h
    port map (
            O => \N__26959\,
            I => \N__26953\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__26956\,
            I => \Inst_core.Inst_sync.filteredInput_7\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__26953\,
            I => \Inst_core.Inst_sync.filteredInput_7\
        );

    \I__5680\ : SRMux
    port map (
            O => \N__26948\,
            I => \N__26945\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__26945\,
            I => \N__26942\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__26942\,
            I => \N__26939\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__26939\,
            I => \Inst_core.Inst_sync.Inst_filter.n4735\
        );

    \I__5676\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26933\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__26933\,
            I => \N__26929\
        );

    \I__5674\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26926\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__26929\,
            I => \N__26923\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__26926\,
            I => \maskRegister_7_adj_1281\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__26923\,
            I => \maskRegister_7_adj_1281\
        );

    \I__5670\ : SRMux
    port map (
            O => \N__26918\,
            I => \N__26915\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__26915\,
            I => \N__26912\
        );

    \I__5668\ : Sp12to4
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__5667\ : Span12Mux_s0_v
    port map (
            O => \N__26909\,
            I => \N__26906\
        );

    \I__5666\ : Odrv12
    port map (
            O => \N__26906\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4752\
        );

    \I__5665\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26899\
        );

    \I__5664\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26896\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__26899\,
            I => \N__26893\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__26896\,
            I => \maskRegister_0_adj_1328\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__26893\,
            I => \maskRegister_0_adj_1328\
        );

    \I__5660\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26884\
        );

    \I__5659\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26881\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__26884\,
            I => \N__26878\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__26881\,
            I => bwd_9
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__26878\,
            I => bwd_9
        );

    \I__5655\ : InMux
    port map (
            O => \N__26873\,
            I => \N__26870\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__26870\,
            I => \Inst_core.Inst_controller.n24\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__26867\,
            I => \Inst_core.Inst_controller.n22_adj_988_cascade_\
        );

    \I__5652\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26861\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__26861\,
            I => \N__26858\
        );

    \I__5650\ : Span4Mux_h
    port map (
            O => \N__26858\,
            I => \N__26853\
        );

    \I__5649\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26848\
        );

    \I__5648\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26848\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__26853\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__26848\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3\
        );

    \I__5645\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26839\
        );

    \I__5644\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26836\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__26839\,
            I => \valueRegister_3_adj_1293\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__26836\,
            I => \valueRegister_3_adj_1293\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__26831\,
            I => \N__26828\
        );

    \I__5640\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26825\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__26822\,
            I => \N__26819\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__5636\ : Odrv4
    port map (
            O => \N__26816\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_3\
        );

    \I__5635\ : SRMux
    port map (
            O => \N__26813\,
            I => \N__26810\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__26810\,
            I => \N__26807\
        );

    \I__5633\ : Span4Mux_h
    port map (
            O => \N__26807\,
            I => \N__26804\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__26804\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4748\
        );

    \I__5631\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26797\
        );

    \I__5630\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26794\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__26797\,
            I => bwd_6
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__26794\,
            I => bwd_6
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__26789\,
            I => \N__26786\
        );

    \I__5626\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26782\
        );

    \I__5625\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26779\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__26782\,
            I => \N__26776\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__26779\,
            I => bwd_5
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__26776\,
            I => bwd_5
        );

    \I__5621\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26768\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__26768\,
            I => \Inst_core.Inst_controller.n23\
        );

    \I__5619\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26761\
        );

    \I__5618\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26758\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__26761\,
            I => bwd_3
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__26758\,
            I => bwd_3
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__26753\,
            I => \N__26749\
        );

    \I__5614\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26746\
        );

    \I__5613\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26743\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__26746\,
            I => bwd_4
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__26743\,
            I => bwd_4
        );

    \I__5610\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26735\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__26735\,
            I => \Inst_core.Inst_controller.n21_adj_989\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__26732\,
            I => \N__26722\
        );

    \I__5607\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26717\
        );

    \I__5606\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26713\
        );

    \I__5605\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26702\
        );

    \I__5604\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26702\
        );

    \I__5603\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26702\
        );

    \I__5602\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26702\
        );

    \I__5601\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26699\
        );

    \I__5600\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26691\
        );

    \I__5599\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26691\
        );

    \I__5598\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26691\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26688\
        );

    \I__5596\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26685\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__26713\,
            I => \N__26682\
        );

    \I__5594\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26677\
        );

    \I__5593\ : InMux
    port map (
            O => \N__26711\,
            I => \N__26677\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__26702\,
            I => \N__26674\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26671\
        );

    \I__5590\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26668\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__26691\,
            I => \N__26665\
        );

    \I__5588\ : Span4Mux_h
    port map (
            O => \N__26688\,
            I => \N__26660\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__26685\,
            I => \N__26660\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__26682\,
            I => \N__26655\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26655\
        );

    \I__5584\ : Span4Mux_v
    port map (
            O => \N__26674\,
            I => \N__26649\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__26671\,
            I => \N__26646\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__26668\,
            I => \N__26643\
        );

    \I__5581\ : Span4Mux_s2_v
    port map (
            O => \N__26665\,
            I => \N__26636\
        );

    \I__5580\ : Span4Mux_v
    port map (
            O => \N__26660\,
            I => \N__26636\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__26655\,
            I => \N__26636\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26633\
        );

    \I__5577\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26630\
        );

    \I__5576\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26627\
        );

    \I__5575\ : Odrv4
    port map (
            O => \N__26649\,
            I => cmd_11
        );

    \I__5574\ : Odrv4
    port map (
            O => \N__26646\,
            I => cmd_11
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__26643\,
            I => cmd_11
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__26636\,
            I => cmd_11
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__26633\,
            I => cmd_11
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__26630\,
            I => cmd_11
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__26627\,
            I => cmd_11
        );

    \I__5568\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26608\
        );

    \I__5567\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26605\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__26608\,
            I => \N__26602\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__26605\,
            I => \configRegister_16_adj_1304\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__26602\,
            I => \configRegister_16_adj_1304\
        );

    \I__5563\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26591\
        );

    \I__5562\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26588\
        );

    \I__5561\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26579\
        );

    \I__5560\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26579\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26576\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__26588\,
            I => \N__26573\
        );

    \I__5557\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26570\
        );

    \I__5556\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26567\
        );

    \I__5555\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26564\
        );

    \I__5554\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26561\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__26579\,
            I => \N__26556\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__26576\,
            I => \N__26556\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__26573\,
            I => \N__26553\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__26570\,
            I => cmd_17
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__26567\,
            I => cmd_17
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__26564\,
            I => cmd_17
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__26561\,
            I => cmd_17
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__26556\,
            I => cmd_17
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__26553\,
            I => cmd_17
        );

    \I__5544\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26531\
        );

    \I__5542\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26528\
        );

    \I__5541\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26525\
        );

    \I__5540\ : CascadeMux
    port map (
            O => \N__26534\,
            I => \N__26521\
        );

    \I__5539\ : Span4Mux_h
    port map (
            O => \N__26531\,
            I => \N__26515\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__26528\,
            I => \N__26512\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__26525\,
            I => \N__26509\
        );

    \I__5536\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26504\
        );

    \I__5535\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26504\
        );

    \I__5534\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26497\
        );

    \I__5533\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26497\
        );

    \I__5532\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26497\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__26515\,
            I => cmd_28
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__26512\,
            I => cmd_28
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__26509\,
            I => cmd_28
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__26504\,
            I => cmd_28
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__26497\,
            I => cmd_28
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__26486\,
            I => \N__26482\
        );

    \I__5525\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26479\
        );

    \I__5524\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26476\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__26479\,
            I => fwd_3
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__26476\,
            I => fwd_3
        );

    \I__5521\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26467\
        );

    \I__5520\ : InMux
    port map (
            O => \N__26470\,
            I => \N__26464\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__26467\,
            I => \N__26461\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__26464\,
            I => \maskRegister_7_adj_1321\
        );

    \I__5517\ : Odrv12
    port map (
            O => \N__26461\,
            I => \maskRegister_7_adj_1321\
        );

    \I__5516\ : SRMux
    port map (
            O => \N__26456\,
            I => \N__26453\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__26453\,
            I => \N__26450\
        );

    \I__5514\ : Span4Mux_h
    port map (
            O => \N__26450\,
            I => \N__26447\
        );

    \I__5513\ : Span4Mux_v
    port map (
            O => \N__26447\,
            I => \N__26444\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__26444\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4759\
        );

    \I__5511\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26438\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26434\
        );

    \I__5509\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26431\
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__26434\,
            I => \maskRegister_0_adj_1368\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__26431\,
            I => \maskRegister_0_adj_1368\
        );

    \I__5506\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26422\
        );

    \I__5505\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26419\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__26422\,
            I => \maskRegister_1_adj_1367\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__26419\,
            I => \maskRegister_1_adj_1367\
        );

    \I__5502\ : InMux
    port map (
            O => \N__26414\,
            I => \N__26410\
        );

    \I__5501\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26407\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__26410\,
            I => \maskRegister_2_adj_1366\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__26407\,
            I => \maskRegister_2_adj_1366\
        );

    \I__5498\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__26399\,
            I => \N__26396\
        );

    \I__5496\ : Span4Mux_v
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__26393\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7_adj_996\
        );

    \I__5494\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26363\
        );

    \I__5493\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26363\
        );

    \I__5492\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26363\
        );

    \I__5491\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26363\
        );

    \I__5490\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26363\
        );

    \I__5489\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26363\
        );

    \I__5488\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26363\
        );

    \I__5487\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26363\
        );

    \I__5486\ : InMux
    port map (
            O => \N__26382\,
            I => \N__26346\
        );

    \I__5485\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26343\
        );

    \I__5484\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26332\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__26363\,
            I => \N__26329\
        );

    \I__5482\ : InMux
    port map (
            O => \N__26362\,
            I => \N__26326\
        );

    \I__5481\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26315\
        );

    \I__5480\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26315\
        );

    \I__5479\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26315\
        );

    \I__5478\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26315\
        );

    \I__5477\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26315\
        );

    \I__5476\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26298\
        );

    \I__5475\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26298\
        );

    \I__5474\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26298\
        );

    \I__5473\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26298\
        );

    \I__5472\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26298\
        );

    \I__5471\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26298\
        );

    \I__5470\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26298\
        );

    \I__5469\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26298\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26295\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__26343\,
            I => \N__26292\
        );

    \I__5466\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26274\
        );

    \I__5465\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26274\
        );

    \I__5464\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26274\
        );

    \I__5463\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26274\
        );

    \I__5462\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26274\
        );

    \I__5461\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26274\
        );

    \I__5460\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26274\
        );

    \I__5459\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26274\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__26332\,
            I => \N__26271\
        );

    \I__5457\ : Span4Mux_s2_v
    port map (
            O => \N__26329\,
            I => \N__26256\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__26326\,
            I => \N__26256\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__26315\,
            I => \N__26256\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__26298\,
            I => \N__26253\
        );

    \I__5453\ : Span4Mux_v
    port map (
            O => \N__26295\,
            I => \N__26248\
        );

    \I__5452\ : Span4Mux_v
    port map (
            O => \N__26292\,
            I => \N__26248\
        );

    \I__5451\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26245\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__26274\,
            I => \N__26241\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__26271\,
            I => \N__26238\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26221\
        );

    \I__5447\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26221\
        );

    \I__5446\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26221\
        );

    \I__5445\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26221\
        );

    \I__5444\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26221\
        );

    \I__5443\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26221\
        );

    \I__5442\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26221\
        );

    \I__5441\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26221\
        );

    \I__5440\ : Span4Mux_v
    port map (
            O => \N__26256\,
            I => \N__26218\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__26253\,
            I => \N__26211\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__26248\,
            I => \N__26211\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__26245\,
            I => \N__26211\
        );

    \I__5436\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26208\
        );

    \I__5435\ : Span4Mux_h
    port map (
            O => \N__26241\,
            I => \N__26203\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__26238\,
            I => \N__26203\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__26221\,
            I => \N__26198\
        );

    \I__5432\ : Span4Mux_h
    port map (
            O => \N__26218\,
            I => \N__26198\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__26211\,
            I => \flagDemux\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__26208\,
            I => \flagDemux\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__26203\,
            I => \flagDemux\
        );

    \I__5428\ : Odrv4
    port map (
            O => \N__26198\,
            I => \flagDemux\
        );

    \I__5427\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26183\
        );

    \I__5426\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26183\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26180\
        );

    \I__5424\ : Odrv12
    port map (
            O => \N__26180\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register\
        );

    \I__5423\ : InMux
    port map (
            O => \N__26177\,
            I => \N__26174\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__26174\,
            I => \N__26170\
        );

    \I__5421\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26167\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__26170\,
            I => \valueRegister_5_adj_1371\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__26167\,
            I => \valueRegister_5_adj_1371\
        );

    \I__5418\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26159\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__26159\,
            I => \N__26156\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__26156\,
            I => \N__26152\
        );

    \I__5415\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26149\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__26152\,
            I => \configRegister_13_adj_1387\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__26149\,
            I => \configRegister_13_adj_1387\
        );

    \I__5412\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26138\
        );

    \I__5411\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26138\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__26138\,
            I => \N__26131\
        );

    \I__5409\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26128\
        );

    \I__5408\ : InMux
    port map (
            O => \N__26136\,
            I => \N__26124\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__26135\,
            I => \N__26121\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__26134\,
            I => \N__26115\
        );

    \I__5405\ : Span4Mux_v
    port map (
            O => \N__26131\,
            I => \N__26107\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__26128\,
            I => \N__26107\
        );

    \I__5403\ : InMux
    port map (
            O => \N__26127\,
            I => \N__26103\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__26124\,
            I => \N__26097\
        );

    \I__5401\ : InMux
    port map (
            O => \N__26121\,
            I => \N__26092\
        );

    \I__5400\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26092\
        );

    \I__5399\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26089\
        );

    \I__5398\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26077\
        );

    \I__5397\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26077\
        );

    \I__5396\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26077\
        );

    \I__5395\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26077\
        );

    \I__5394\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26072\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__26107\,
            I => \N__26069\
        );

    \I__5392\ : InMux
    port map (
            O => \N__26106\,
            I => \N__26066\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__26103\,
            I => \N__26063\
        );

    \I__5390\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26060\
        );

    \I__5389\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26055\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26100\,
            I => \N__26055\
        );

    \I__5387\ : Span4Mux_v
    port map (
            O => \N__26097\,
            I => \N__26050\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__26092\,
            I => \N__26050\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__26089\,
            I => \N__26045\
        );

    \I__5384\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26038\
        );

    \I__5383\ : InMux
    port map (
            O => \N__26087\,
            I => \N__26038\
        );

    \I__5382\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26038\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__26077\,
            I => \N__26035\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26030\
        );

    \I__5379\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26030\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__26072\,
            I => \N__26027\
        );

    \I__5377\ : Sp12to4
    port map (
            O => \N__26069\,
            I => \N__26021\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26066\,
            I => \N__26021\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__26063\,
            I => \N__26012\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__26060\,
            I => \N__26012\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__26055\,
            I => \N__26012\
        );

    \I__5372\ : Span4Mux_h
    port map (
            O => \N__26050\,
            I => \N__26012\
        );

    \I__5371\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26007\
        );

    \I__5370\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26007\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__26045\,
            I => \N__26000\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__26038\,
            I => \N__26000\
        );

    \I__5367\ : Span4Mux_s1_v
    port map (
            O => \N__26035\,
            I => \N__26000\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26030\,
            I => \N__25995\
        );

    \I__5365\ : Span4Mux_v
    port map (
            O => \N__26027\,
            I => \N__25995\
        );

    \I__5364\ : InMux
    port map (
            O => \N__26026\,
            I => \N__25992\
        );

    \I__5363\ : Span12Mux_s8_h
    port map (
            O => \N__26021\,
            I => \N__25989\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__26012\,
            I => \N__25986\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__26007\,
            I => \N__25979\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__26000\,
            I => \N__25979\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__25995\,
            I => \N__25979\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__25992\,
            I => wrtrigcfg_3
        );

    \I__5357\ : Odrv12
    port map (
            O => \N__25989\,
            I => wrtrigcfg_3
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__25986\,
            I => wrtrigcfg_3
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__25979\,
            I => wrtrigcfg_3
        );

    \I__5354\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25966\
        );

    \I__5353\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25963\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__25966\,
            I => \N__25960\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__25963\,
            I => \configRegister_16_adj_1384\
        );

    \I__5350\ : Odrv4
    port map (
            O => \N__25960\,
            I => \configRegister_16_adj_1384\
        );

    \I__5349\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25952\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__25952\,
            I => \N__25948\
        );

    \I__5347\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25945\
        );

    \I__5346\ : Odrv4
    port map (
            O => \N__25948\,
            I => \configRegister_12_adj_1348\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__25945\,
            I => \configRegister_12_adj_1348\
        );

    \I__5344\ : SRMux
    port map (
            O => \N__25940\,
            I => \N__25929\
        );

    \I__5343\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25920\
        );

    \I__5342\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25920\
        );

    \I__5341\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25920\
        );

    \I__5340\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25920\
        );

    \I__5339\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25911\
        );

    \I__5338\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25911\
        );

    \I__5337\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25911\
        );

    \I__5336\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25911\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__25929\,
            I => \N__25908\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__25920\,
            I => \N__25903\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__25911\,
            I => \N__25903\
        );

    \I__5332\ : Span12Mux_s11_v
    port map (
            O => \N__25908\,
            I => \N__25898\
        );

    \I__5331\ : Span12Mux_s4_v
    port map (
            O => \N__25903\,
            I => \N__25898\
        );

    \I__5330\ : Odrv12
    port map (
            O => \N__25898\,
            I => \Inst_core.arm\
        );

    \I__5329\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25891\
        );

    \I__5328\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25888\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__25891\,
            I => \maskRegister_5_adj_1323\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__25888\,
            I => \maskRegister_5_adj_1323\
        );

    \I__5325\ : SRMux
    port map (
            O => \N__25883\,
            I => \N__25880\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__25880\,
            I => \N__25877\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__25874\,
            I => \N__25871\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__25871\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4757\
        );

    \I__5320\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25864\
        );

    \I__5319\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25861\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__25864\,
            I => \maskRegister_6_adj_1322\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__25861\,
            I => \maskRegister_6_adj_1322\
        );

    \I__5316\ : CascadeMux
    port map (
            O => \N__25856\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n2_cascade_\
        );

    \I__5315\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25850\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__25850\,
            I => \N__25847\
        );

    \I__5313\ : Span4Mux_v
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__25844\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register\
        );

    \I__5311\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25835\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__25835\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n100\
        );

    \I__5308\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25828\
        );

    \I__5307\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25825\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__25828\,
            I => \N__25822\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__25825\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n553\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__25822\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n553\
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__25817\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n100_cascade_\
        );

    \I__5302\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__25811\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__25808\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n2_cascade_\
        );

    \I__5299\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25798\
        );

    \I__5297\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25795\
        );

    \I__5296\ : Span4Mux_s3_h
    port map (
            O => \N__25798\,
            I => \N__25792\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__25795\,
            I => \configRegister_17_adj_1383\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__25792\,
            I => \configRegister_17_adj_1383\
        );

    \I__5293\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25784\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__25781\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n100\
        );

    \I__5290\ : CascadeMux
    port map (
            O => \N__25778\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n100_cascade_\
        );

    \I__5289\ : CascadeMux
    port map (
            O => \N__25775\,
            I => \N__25771\
        );

    \I__5288\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25768\
        );

    \I__5287\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25762\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__25765\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n759\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__25762\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n759\
        );

    \I__5283\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__25751\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n770\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__25748\,
            I => \N__25740\
        );

    \I__5279\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25736\
        );

    \I__5278\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25727\
        );

    \I__5277\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25727\
        );

    \I__5276\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25727\
        );

    \I__5275\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25727\
        );

    \I__5274\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25722\
        );

    \I__5273\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25722\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25719\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__25727\,
            I => \N__25716\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__25722\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.state_1\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__25719\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.state_1\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__25716\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.state_1\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__25709\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n770_cascade_\
        );

    \I__5266\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25703\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__5264\ : Odrv12
    port map (
            O => \N__25700\,
            I => \Inst_core.n6713\
        );

    \I__5263\ : CEMux
    port map (
            O => \N__25697\,
            I => \N__25693\
        );

    \I__5262\ : CEMux
    port map (
            O => \N__25696\,
            I => \N__25690\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__25693\,
            I => \N__25687\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__25690\,
            I => \N__25684\
        );

    \I__5259\ : Span4Mux_v
    port map (
            O => \N__25687\,
            I => \N__25681\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__25684\,
            I => \N__25678\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__25681\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4076\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__25678\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4076\
        );

    \I__5255\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25669\
        );

    \I__5254\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25666\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25663\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__25666\,
            I => \configRegister_17_adj_1303\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__25663\,
            I => \configRegister_17_adj_1303\
        );

    \I__5250\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25655\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__25655\,
            I => \N__25652\
        );

    \I__5248\ : Span4Mux_s2_v
    port map (
            O => \N__25652\,
            I => \N__25648\
        );

    \I__5247\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25645\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__25648\,
            I => \configRegister_4_adj_1356\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__25645\,
            I => \configRegister_4_adj_1356\
        );

    \I__5244\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25636\
        );

    \I__5243\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25633\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25630\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__25633\,
            I => \maskRegister_5_adj_1363\
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__25630\,
            I => \maskRegister_5_adj_1363\
        );

    \I__5239\ : SRMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__25622\,
            I => \N__25619\
        );

    \I__5237\ : Span4Mux_v
    port map (
            O => \N__25619\,
            I => \N__25616\
        );

    \I__5236\ : Odrv4
    port map (
            O => \N__25616\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4764\
        );

    \I__5235\ : CascadeMux
    port map (
            O => \N__25613\,
            I => \N__25610\
        );

    \I__5234\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25605\
        );

    \I__5233\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25600\
        );

    \I__5232\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25600\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__25605\,
            I => \N__25594\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__25600\,
            I => \N__25594\
        );

    \I__5229\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25590\
        );

    \I__5228\ : Span4Mux_v
    port map (
            O => \N__25594\,
            I => \N__25584\
        );

    \I__5227\ : InMux
    port map (
            O => \N__25593\,
            I => \N__25581\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__25590\,
            I => \N__25578\
        );

    \I__5225\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25571\
        );

    \I__5224\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25571\
        );

    \I__5223\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25571\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__25584\,
            I => cmd_18
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__25581\,
            I => cmd_18
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__25578\,
            I => cmd_18
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__25571\,
            I => cmd_18
        );

    \I__5218\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__25559\,
            I => \N__25555\
        );

    \I__5216\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25552\
        );

    \I__5215\ : Odrv4
    port map (
            O => \N__25555\,
            I => \configRegister_13_adj_1347\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__25552\,
            I => \configRegister_13_adj_1347\
        );

    \I__5213\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25544\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__25544\,
            I => \N__25540\
        );

    \I__5211\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25537\
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__25540\,
            I => \configRegister_14_adj_1386\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__25537\,
            I => \configRegister_14_adj_1386\
        );

    \I__5208\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25529\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__25529\,
            I => \N__25524\
        );

    \I__5206\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25519\
        );

    \I__5205\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25519\
        );

    \I__5204\ : Odrv4
    port map (
            O => \N__25524\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__25519\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__25514\,
            I => \N__25508\
        );

    \I__5201\ : InMux
    port map (
            O => \N__25513\,
            I => \N__25504\
        );

    \I__5200\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25501\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__25511\,
            I => \N__25497\
        );

    \I__5198\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25494\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__25507\,
            I => \N__25491\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__25504\,
            I => \N__25483\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__25501\,
            I => \N__25483\
        );

    \I__5194\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25480\
        );

    \I__5193\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25477\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__25494\,
            I => \N__25474\
        );

    \I__5191\ : InMux
    port map (
            O => \N__25491\,
            I => \N__25471\
        );

    \I__5190\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25468\
        );

    \I__5189\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25465\
        );

    \I__5188\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25462\
        );

    \I__5187\ : Span4Mux_v
    port map (
            O => \N__25483\,
            I => \N__25459\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25456\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__25477\,
            I => \N__25452\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__25474\,
            I => \N__25449\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__25471\,
            I => \N__25446\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__25468\,
            I => \N__25441\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__25465\,
            I => \N__25441\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__25462\,
            I => \N__25438\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__25459\,
            I => \N__25433\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__25456\,
            I => \N__25433\
        );

    \I__5177\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25430\
        );

    \I__5176\ : Span4Mux_v
    port map (
            O => \N__25452\,
            I => \N__25425\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__25449\,
            I => \N__25425\
        );

    \I__5174\ : Span12Mux_v
    port map (
            O => \N__25446\,
            I => \N__25422\
        );

    \I__5173\ : Span12Mux_v
    port map (
            O => \N__25441\,
            I => \N__25419\
        );

    \I__5172\ : Span4Mux_v
    port map (
            O => \N__25438\,
            I => \N__25414\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__25433\,
            I => \N__25414\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__25430\,
            I => \memoryOut_5\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__25425\,
            I => \memoryOut_5\
        );

    \I__5168\ : Odrv12
    port map (
            O => \N__25422\,
            I => \memoryOut_5\
        );

    \I__5167\ : Odrv12
    port map (
            O => \N__25419\,
            I => \memoryOut_5\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__25414\,
            I => \memoryOut_5\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__5164\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25394\
        );

    \I__5163\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25394\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__25394\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n554\
        );

    \I__5161\ : CascadeMux
    port map (
            O => \N__25391\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n22_cascade_\
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__25388\,
            I => \Inst_core.n8515_cascade_\
        );

    \I__5159\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25379\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25379\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__25379\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n451\
        );

    \I__5156\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25370\
        );

    \I__5155\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25370\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__25370\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n760\
        );

    \I__5153\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25358\
        );

    \I__5152\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25349\
        );

    \I__5151\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25349\
        );

    \I__5150\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25349\
        );

    \I__5149\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25349\
        );

    \I__5148\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25344\
        );

    \I__5147\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25344\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25341\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__25349\,
            I => \N__25338\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__25344\,
            I => \N__25331\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__25341\,
            I => \N__25331\
        );

    \I__5142\ : Span4Mux_s2_v
    port map (
            O => \N__25338\,
            I => \N__25331\
        );

    \I__5141\ : Odrv4
    port map (
            O => \N__25331\,
            I => \Inst_core.n31\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__25328\,
            I => \N__25317\
        );

    \I__5139\ : CascadeMux
    port map (
            O => \N__25327\,
            I => \N__25313\
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__25326\,
            I => \N__25309\
        );

    \I__5137\ : CascadeMux
    port map (
            O => \N__25325\,
            I => \N__25305\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__25324\,
            I => \N__25302\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__25323\,
            I => \N__25298\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__25322\,
            I => \N__25294\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__25321\,
            I => \N__25290\
        );

    \I__5132\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25273\
        );

    \I__5131\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25273\
        );

    \I__5130\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25273\
        );

    \I__5129\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25273\
        );

    \I__5128\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25273\
        );

    \I__5127\ : InMux
    port map (
            O => \N__25309\,
            I => \N__25273\
        );

    \I__5126\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25273\
        );

    \I__5125\ : InMux
    port map (
            O => \N__25305\,
            I => \N__25273\
        );

    \I__5124\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25258\
        );

    \I__5123\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25258\
        );

    \I__5122\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25258\
        );

    \I__5121\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25258\
        );

    \I__5120\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25258\
        );

    \I__5119\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25258\
        );

    \I__5118\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25258\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__25273\,
            I => \N__25255\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25252\
        );

    \I__5115\ : Span4Mux_h
    port map (
            O => \N__25255\,
            I => \N__25249\
        );

    \I__5114\ : Span4Mux_h
    port map (
            O => \N__25252\,
            I => \N__25246\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__25249\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n1765\
        );

    \I__5112\ : Odrv4
    port map (
            O => \N__25246\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n1765\
        );

    \I__5111\ : InMux
    port map (
            O => \N__25241\,
            I => \N__25238\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__25238\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n667\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__25235\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n667_cascade_\
        );

    \I__5108\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__25229\,
            I => \N__25222\
        );

    \I__5106\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25213\
        );

    \I__5105\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25213\
        );

    \I__5104\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25213\
        );

    \I__5103\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25213\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__25222\,
            I => \Inst_core.n31_adj_1174\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__25213\,
            I => \Inst_core.n31_adj_1174\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__25208\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n100_cascade_\
        );

    \I__5099\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25199\
        );

    \I__5098\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25199\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__25199\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n656\
        );

    \I__5096\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25193\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__25193\,
            I => \Inst_core.n8518\
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__5093\ : InMux
    port map (
            O => \N__25187\,
            I => \N__25179\
        );

    \I__5092\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25176\
        );

    \I__5091\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25173\
        );

    \I__5090\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25170\
        );

    \I__5089\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25165\
        );

    \I__5088\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25165\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__25179\,
            I => \Inst_core.state_1_adj_1134\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__25176\,
            I => \Inst_core.state_1_adj_1134\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__25173\,
            I => \Inst_core.state_1_adj_1134\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__25170\,
            I => \Inst_core.state_1_adj_1134\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__25165\,
            I => \Inst_core.state_1_adj_1134\
        );

    \I__5082\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25148\
        );

    \I__5081\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25148\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__25148\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n657\
        );

    \I__5079\ : InMux
    port map (
            O => \N__25145\,
            I => \N__25141\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__25144\,
            I => \N__25138\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__25141\,
            I => \N__25134\
        );

    \I__5076\ : InMux
    port map (
            O => \N__25138\,
            I => \N__25129\
        );

    \I__5075\ : InMux
    port map (
            O => \N__25137\,
            I => \N__25129\
        );

    \I__5074\ : Odrv4
    port map (
            O => \N__25134\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__25129\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4\
        );

    \I__5072\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__25121\,
            I => \N__25116\
        );

    \I__5070\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25111\
        );

    \I__5069\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25111\
        );

    \I__5068\ : Odrv4
    port map (
            O => \N__25116\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__25111\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__25106\,
            I => \N__25103\
        );

    \I__5065\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25100\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25097\
        );

    \I__5063\ : Span4Mux_v
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__25094\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_7\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__25091\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n8844_cascade_\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__25085\,
            I => \Inst_core.Inst_decoder.n6\
        );

    \I__5058\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__25073\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9052\
        );

    \I__5054\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25067\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25063\
        );

    \I__5052\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__5051\ : Odrv12
    port map (
            O => \N__25063\,
            I => \valueRegister_1_adj_1335\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__25060\,
            I => \valueRegister_1_adj_1335\
        );

    \I__5049\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25051\
        );

    \I__5048\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25047\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__25051\,
            I => \N__25044\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25050\,
            I => \N__25041\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__25047\,
            I => \N__25036\
        );

    \I__5044\ : Span4Mux_s3_v
    port map (
            O => \N__25044\,
            I => \N__25036\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__25041\,
            I => divider_20
        );

    \I__5042\ : Odrv4
    port map (
            O => \N__25036\,
            I => divider_20
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__25031\,
            I => \N__25028\
        );

    \I__5040\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25024\
        );

    \I__5039\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25020\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__25024\,
            I => \N__25017\
        );

    \I__5037\ : InMux
    port map (
            O => \N__25023\,
            I => \N__25014\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__25020\,
            I => divider_21
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__25017\,
            I => divider_21
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__25014\,
            I => divider_21
        );

    \I__5033\ : InMux
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__25004\,
            I => \N__25001\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__25001\,
            I => \Inst_core.Inst_sampler.n8598\
        );

    \I__5030\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24995\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__24992\,
            I => \Inst_core.Inst_sampler.n8602\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__24989\,
            I => \Inst_core.Inst_sampler.n8600_cascade_\
        );

    \I__5026\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__24983\,
            I => \Inst_core.Inst_sampler.n8604\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__24980\,
            I => \N__24977\
        );

    \I__5023\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__24974\,
            I => \N__24970\
        );

    \I__5021\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24967\
        );

    \I__5020\ : Span4Mux_s3_v
    port map (
            O => \N__24970\,
            I => \N__24964\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__24967\,
            I => \N__24959\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__24964\,
            I => \N__24959\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__24959\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelL16\
        );

    \I__5016\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24953\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__24953\,
            I => \N__24950\
        );

    \I__5014\ : Span12Mux_s6_h
    port map (
            O => \N__24950\,
            I => \N__24946\
        );

    \I__5013\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24943\
        );

    \I__5012\ : Odrv12
    port map (
            O => \N__24946\,
            I => \configRegister_24_adj_1338\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__24943\,
            I => \configRegister_24_adj_1338\
        );

    \I__5010\ : InMux
    port map (
            O => \N__24938\,
            I => \N__24932\
        );

    \I__5009\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24932\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__24932\,
            I => \N__24929\
        );

    \I__5007\ : Span4Mux_h
    port map (
            O => \N__24929\,
            I => \N__24925\
        );

    \I__5006\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__24925\,
            I => \N__24919\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__24922\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16\
        );

    \I__5003\ : Odrv4
    port map (
            O => \N__24919\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16\
        );

    \I__5002\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24909\
        );

    \I__5001\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24904\
        );

    \I__5000\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24904\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__24909\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__24904\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__4996\ : InMux
    port map (
            O => \N__24896\,
            I => \N__24892\
        );

    \I__4995\ : InMux
    port map (
            O => \N__24895\,
            I => \N__24889\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__24892\,
            I => \N__24883\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__24889\,
            I => \N__24883\
        );

    \I__4992\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24880\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__24883\,
            I => \N__24877\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__24880\,
            I => divider_9
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__24877\,
            I => divider_9
        );

    \I__4988\ : CascadeMux
    port map (
            O => \N__24872\,
            I => \N__24868\
        );

    \I__4987\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24864\
        );

    \I__4986\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24861\
        );

    \I__4985\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24858\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24853\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24853\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__24858\,
            I => divider_7
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__24853\,
            I => divider_7
        );

    \I__4980\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__24845\,
            I => \Inst_core.Inst_sampler.n29\
        );

    \I__4978\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__24836\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_7\
        );

    \I__4975\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24830\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__24830\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_4\
        );

    \I__4973\ : InMux
    port map (
            O => \N__24827\,
            I => \N__24824\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__24824\,
            I => \N__24820\
        );

    \I__4971\ : InMux
    port map (
            O => \N__24823\,
            I => \N__24817\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__24820\,
            I => \valueRegister_5_adj_1331\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__24817\,
            I => \valueRegister_5_adj_1331\
        );

    \I__4968\ : CascadeMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__4967\ : InMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__24806\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_5\
        );

    \I__4965\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24798\
        );

    \I__4964\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24795\
        );

    \I__4963\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24792\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__24798\,
            I => divider_15
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__24795\,
            I => divider_15
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__24792\,
            I => divider_15
        );

    \I__4959\ : CascadeMux
    port map (
            O => \N__24785\,
            I => \N__24782\
        );

    \I__4958\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24779\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24775\
        );

    \I__4956\ : CascadeMux
    port map (
            O => \N__24778\,
            I => \N__24772\
        );

    \I__4955\ : Span4Mux_h
    port map (
            O => \N__24775\,
            I => \N__24768\
        );

    \I__4954\ : InMux
    port map (
            O => \N__24772\,
            I => \N__24765\
        );

    \I__4953\ : InMux
    port map (
            O => \N__24771\,
            I => \N__24762\
        );

    \I__4952\ : Span4Mux_v
    port map (
            O => \N__24768\,
            I => \N__24759\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__24765\,
            I => \N__24756\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__24762\,
            I => divider_13
        );

    \I__4949\ : Odrv4
    port map (
            O => \N__24759\,
            I => divider_13
        );

    \I__4948\ : Odrv12
    port map (
            O => \N__24756\,
            I => divider_13
        );

    \I__4947\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24744\
        );

    \I__4946\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24741\
        );

    \I__4945\ : InMux
    port map (
            O => \N__24747\,
            I => \N__24738\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__24744\,
            I => divider_16
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__24741\,
            I => divider_16
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__24738\,
            I => divider_16
        );

    \I__4941\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__24728\,
            I => \Inst_core.Inst_sampler.n32\
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__24725\,
            I => \N__24721\
        );

    \I__4938\ : CascadeMux
    port map (
            O => \N__24724\,
            I => \N__24718\
        );

    \I__4937\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24715\
        );

    \I__4936\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24712\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__24715\,
            I => \N__24706\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__24712\,
            I => \N__24706\
        );

    \I__4933\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24703\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__24706\,
            I => \N__24700\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__24703\,
            I => divider_14
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__24700\,
            I => divider_14
        );

    \I__4929\ : CascadeMux
    port map (
            O => \N__24695\,
            I => \Inst_core.Inst_sampler.n8596_cascade_\
        );

    \I__4928\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__24689\,
            I => \Inst_core.Inst_sampler.n8590\
        );

    \I__4926\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24681\
        );

    \I__4925\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24678\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__24684\,
            I => \N__24675\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__24681\,
            I => \N__24670\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__24678\,
            I => \N__24670\
        );

    \I__4921\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24665\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__24670\,
            I => \N__24659\
        );

    \I__4919\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24654\
        );

    \I__4918\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24654\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__24665\,
            I => \N__24651\
        );

    \I__4916\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24644\
        );

    \I__4915\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24644\
        );

    \I__4914\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24644\
        );

    \I__4913\ : Odrv4
    port map (
            O => \N__24659\,
            I => cmd_29
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__24654\,
            I => cmd_29
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__24651\,
            I => cmd_29
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__24644\,
            I => cmd_29
        );

    \I__4909\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__24632\,
            I => \syncedInput_0\
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__4906\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24623\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__24623\,
            I => \N__24620\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__24617\,
            I => \syncedInput_1\
        );

    \I__4902\ : CascadeMux
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__4901\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24604\
        );

    \I__4899\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24601\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__24604\,
            I => \valueRegister_4_adj_1332\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__24601\,
            I => \valueRegister_4_adj_1332\
        );

    \I__4896\ : SRMux
    port map (
            O => \N__24596\,
            I => \N__24593\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__24593\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4756\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__24590\,
            I => \Inst_core.Inst_sampler.n31_adj_995_cascade_\
        );

    \I__4893\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__4891\ : Span4Mux_h
    port map (
            O => \N__24581\,
            I => \N__24577\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__24580\,
            I => \N__24574\
        );

    \I__4889\ : Span4Mux_v
    port map (
            O => \N__24577\,
            I => \N__24570\
        );

    \I__4888\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24565\
        );

    \I__4887\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24565\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__24570\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__24565\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__4883\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__24554\,
            I => \N__24551\
        );

    \I__4881\ : Span4Mux_h
    port map (
            O => \N__24551\,
            I => \N__24547\
        );

    \I__4880\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24544\
        );

    \I__4879\ : Odrv4
    port map (
            O => \N__24547\,
            I => \valueRegister_4_adj_1292\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__24544\,
            I => \valueRegister_4_adj_1292\
        );

    \I__4877\ : SRMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__4875\ : Span4Mux_v
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__24530\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4749\
        );

    \I__4873\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__24524\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_5\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__4870\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__4868\ : Odrv12
    port map (
            O => \N__24512\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_7\
        );

    \I__4867\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24506\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__24506\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_4\
        );

    \I__4865\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24499\
        );

    \I__4864\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24496\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__24499\,
            I => \N__24493\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__24496\,
            I => fwd_12
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__24493\,
            I => fwd_12
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__24488\,
            I => \N__24485\
        );

    \I__4859\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24481\
        );

    \I__4858\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24475\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__24478\,
            I => fwd_1
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__24475\,
            I => fwd_1
        );

    \I__4854\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__24467\,
            I => \Inst_core.Inst_controller.n13\
        );

    \I__4852\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24460\
        );

    \I__4851\ : InMux
    port map (
            O => \N__24463\,
            I => \N__24457\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__24460\,
            I => \N__24454\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__24457\,
            I => bwd_10
        );

    \I__4848\ : Odrv12
    port map (
            O => \N__24454\,
            I => bwd_10
        );

    \I__4847\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__24446\,
            I => \Inst_core.Inst_controller.n14\
        );

    \I__4845\ : InMux
    port map (
            O => \N__24443\,
            I => \N__24440\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__4843\ : Span4Mux_v
    port map (
            O => \N__24437\,
            I => \N__24433\
        );

    \I__4842\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24430\
        );

    \I__4841\ : Sp12to4
    port map (
            O => \N__24433\,
            I => \N__24427\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__24430\,
            I => fwd_8
        );

    \I__4839\ : Odrv12
    port map (
            O => \N__24427\,
            I => fwd_8
        );

    \I__4838\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24419\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__24419\,
            I => \Inst_core.Inst_controller.n11\
        );

    \I__4836\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24413\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__4834\ : Span4Mux_h
    port map (
            O => \N__24410\,
            I => \N__24407\
        );

    \I__4833\ : Span4Mux_h
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__24404\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n14\
        );

    \I__4831\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__24398\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n11\
        );

    \I__4829\ : CascadeMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__4828\ : InMux
    port map (
            O => \N__24392\,
            I => \N__24385\
        );

    \I__4827\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24385\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__24390\,
            I => \N__24382\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__24385\,
            I => \N__24379\
        );

    \I__4824\ : InMux
    port map (
            O => \N__24382\,
            I => \N__24376\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__24379\,
            I => cmd_37
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__24376\,
            I => cmd_37
        );

    \I__4821\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24368\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__24368\,
            I => \N__24363\
        );

    \I__4819\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24358\
        );

    \I__4818\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24358\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__24363\,
            I => cmd_36
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__24358\,
            I => cmd_36
        );

    \I__4815\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24350\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__24350\,
            I => \N__24347\
        );

    \I__4813\ : Span12Mux_s3_v
    port map (
            O => \N__24347\,
            I => \N__24343\
        );

    \I__4812\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24340\
        );

    \I__4811\ : Odrv12
    port map (
            O => \N__24343\,
            I => \configRegister_6_adj_1354\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__24340\,
            I => \configRegister_6_adj_1354\
        );

    \I__4809\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__24329\,
            I => \N__24325\
        );

    \I__4806\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24322\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__24325\,
            I => \valueRegister_5_adj_1291\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__24322\,
            I => \valueRegister_5_adj_1291\
        );

    \I__4803\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24314\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__4801\ : Span4Mux_h
    port map (
            O => \N__24311\,
            I => \N__24306\
        );

    \I__4800\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24301\
        );

    \I__4799\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24301\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__24306\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__24301\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5\
        );

    \I__4796\ : SRMux
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__24293\,
            I => \N__24290\
        );

    \I__4794\ : Span4Mux_h
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__24287\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4750\
        );

    \I__4792\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24280\
        );

    \I__4791\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24277\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__24280\,
            I => \N__24274\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__24277\,
            I => bwd_11
        );

    \I__4788\ : Odrv12
    port map (
            O => \N__24274\,
            I => bwd_11
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__24269\,
            I => \N__24266\
        );

    \I__4786\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24262\
        );

    \I__4785\ : InMux
    port map (
            O => \N__24265\,
            I => \N__24259\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__24262\,
            I => \N__24256\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__24259\,
            I => bwd_8
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__24256\,
            I => bwd_8
        );

    \I__4781\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24247\
        );

    \I__4780\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24244\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__24247\,
            I => fwd_11
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__24244\,
            I => fwd_11
        );

    \I__4777\ : CascadeMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__4776\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24232\
        );

    \I__4775\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24229\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24224\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24224\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__24224\,
            I => fwd_4
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__24221\,
            I => \Inst_core.Inst_controller.n18_cascade_\
        );

    \I__4770\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24215\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__24215\,
            I => \Inst_core.Inst_controller.n21\
        );

    \I__4768\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24208\
        );

    \I__4767\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24205\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__24208\,
            I => fwd_13
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__24205\,
            I => fwd_13
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__24200\,
            I => \N__24196\
        );

    \I__4763\ : InMux
    port map (
            O => \N__24199\,
            I => \N__24193\
        );

    \I__4762\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24190\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__24193\,
            I => fwd_9
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__24190\,
            I => fwd_9
        );

    \I__4759\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24182\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__24182\,
            I => \Inst_core.Inst_controller.n15\
        );

    \I__4757\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24172\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__24178\,
            I => \N__24169\
        );

    \I__4755\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24163\
        );

    \I__4754\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24163\
        );

    \I__4753\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24160\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__24172\,
            I => \N__24157\
        );

    \I__4751\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24154\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__24168\,
            I => \N__24149\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__24163\,
            I => \N__24146\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__24160\,
            I => \N__24143\
        );

    \I__4747\ : Span4Mux_v
    port map (
            O => \N__24157\,
            I => \N__24138\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24138\
        );

    \I__4745\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24135\
        );

    \I__4744\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24130\
        );

    \I__4743\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24130\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__24146\,
            I => cmd_30
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__24143\,
            I => cmd_30
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__24138\,
            I => cmd_30
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__24135\,
            I => cmd_30
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__24130\,
            I => cmd_30
        );

    \I__4737\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24112\
        );

    \I__4736\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24112\
        );

    \I__4735\ : InMux
    port map (
            O => \N__24117\,
            I => \N__24109\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__24112\,
            I => \N__24106\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__24109\,
            I => \configRegister_22\
        );

    \I__4732\ : Odrv12
    port map (
            O => \N__24106\,
            I => \configRegister_22\
        );

    \I__4731\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24096\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24093\
        );

    \I__4729\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24090\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__24096\,
            I => cmd_33
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__24093\,
            I => cmd_33
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__24090\,
            I => cmd_33
        );

    \I__4725\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24080\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__24080\,
            I => \N__24077\
        );

    \I__4723\ : Span4Mux_v
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__24074\,
            I => \N__24070\
        );

    \I__4721\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24067\
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__24070\,
            I => \configRegister_9_adj_1391\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__24067\,
            I => \configRegister_9_adj_1391\
        );

    \I__4718\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24058\
        );

    \I__4717\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24055\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__24058\,
            I => \N__24050\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__24055\,
            I => \N__24050\
        );

    \I__4714\ : Span4Mux_v
    port map (
            O => \N__24050\,
            I => \N__24046\
        );

    \I__4713\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24043\
        );

    \I__4712\ : Span4Mux_h
    port map (
            O => \N__24046\,
            I => \N__24040\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__24043\,
            I => cmd_38
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__24040\,
            I => cmd_38
        );

    \I__4709\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24031\
        );

    \I__4708\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24028\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__24031\,
            I => \N__24025\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__24028\,
            I => \N__24020\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__24025\,
            I => \N__24020\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__24020\,
            I => \Inst_core.Inst_controller.fwd_14\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24014\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__4701\ : Span4Mux_s2_v
    port map (
            O => \N__24011\,
            I => \N__24007\
        );

    \I__4700\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24004\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__24007\,
            I => \configRegister_8_adj_1352\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__24004\,
            I => \configRegister_8_adj_1352\
        );

    \I__4697\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23994\
        );

    \I__4696\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23989\
        );

    \I__4695\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23986\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__23994\,
            I => \N__23982\
        );

    \I__4693\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23979\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__23992\,
            I => \N__23975\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23971\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__23986\,
            I => \N__23968\
        );

    \I__4689\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23965\
        );

    \I__4688\ : Span4Mux_v
    port map (
            O => \N__23982\,
            I => \N__23960\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__23979\,
            I => \N__23960\
        );

    \I__4686\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23957\
        );

    \I__4685\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23952\
        );

    \I__4684\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23952\
        );

    \I__4683\ : Odrv12
    port map (
            O => \N__23971\,
            I => cmd_16
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__23968\,
            I => cmd_16
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__23965\,
            I => cmd_16
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__23960\,
            I => cmd_16
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__23957\,
            I => cmd_16
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__23952\,
            I => cmd_16
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__4676\ : InMux
    port map (
            O => \N__23936\,
            I => \N__23933\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__23933\,
            I => \N__23929\
        );

    \I__4674\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23926\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__23929\,
            I => \configRegister_15_adj_1345\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__23926\,
            I => \configRegister_15_adj_1345\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__23921\,
            I => \N__23913\
        );

    \I__4670\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23904\
        );

    \I__4669\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23904\
        );

    \I__4668\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23904\
        );

    \I__4667\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23901\
        );

    \I__4666\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23892\
        );

    \I__4665\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23892\
        );

    \I__4664\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23892\
        );

    \I__4663\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23892\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__23904\,
            I => \N__23885\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__23901\,
            I => \N__23885\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__23892\,
            I => \N__23885\
        );

    \I__4659\ : Odrv12
    port map (
            O => \N__23885\,
            I => wrtrigmask_3
        );

    \I__4658\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23875\
        );

    \I__4656\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23872\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__23875\,
            I => \configRegister_12_adj_1388\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__23872\,
            I => \configRegister_12_adj_1388\
        );

    \I__4653\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__23864\,
            I => \N__23860\
        );

    \I__4651\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__23860\,
            I => \configRegister_5_adj_1355\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__23857\,
            I => \configRegister_5_adj_1355\
        );

    \I__4648\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23849\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__23849\,
            I => \N__23845\
        );

    \I__4646\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23842\
        );

    \I__4645\ : Odrv12
    port map (
            O => \N__23845\,
            I => \configRegister_14_adj_1346\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__23842\,
            I => \configRegister_14_adj_1346\
        );

    \I__4643\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23834\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23830\
        );

    \I__4641\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23827\
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__23830\,
            I => \configRegister_9_adj_1351\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__23827\,
            I => \configRegister_9_adj_1351\
        );

    \I__4638\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23818\
        );

    \I__4637\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23815\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__23818\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__23815\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12\
        );

    \I__4634\ : InMux
    port map (
            O => \N__23810\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7910\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__23807\,
            I => \N__23804\
        );

    \I__4632\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23800\
        );

    \I__4631\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23797\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__23800\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__23797\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13\
        );

    \I__4628\ : InMux
    port map (
            O => \N__23792\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7911\
        );

    \I__4627\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23785\
        );

    \I__4626\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23782\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__23785\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__23782\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14\
        );

    \I__4623\ : InMux
    port map (
            O => \N__23777\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7912\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__23774\,
            I => \N__23766\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__23773\,
            I => \N__23762\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__23772\,
            I => \N__23758\
        );

    \I__4619\ : CascadeMux
    port map (
            O => \N__23771\,
            I => \N__23754\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__23770\,
            I => \N__23748\
        );

    \I__4617\ : InMux
    port map (
            O => \N__23769\,
            I => \N__23745\
        );

    \I__4616\ : InMux
    port map (
            O => \N__23766\,
            I => \N__23730\
        );

    \I__4615\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23730\
        );

    \I__4614\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23730\
        );

    \I__4613\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23730\
        );

    \I__4612\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23730\
        );

    \I__4611\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23730\
        );

    \I__4610\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23730\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__23753\,
            I => \N__23726\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__23752\,
            I => \N__23722\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__23751\,
            I => \N__23718\
        );

    \I__4606\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23715\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__23745\,
            I => \N__23710\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23710\
        );

    \I__4603\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23697\
        );

    \I__4602\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23697\
        );

    \I__4601\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23697\
        );

    \I__4600\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23697\
        );

    \I__4599\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23697\
        );

    \I__4598\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23697\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23694\
        );

    \I__4596\ : Odrv4
    port map (
            O => \N__23710\,
            I => \Inst_core.n1639\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__23697\,
            I => \Inst_core.n1639\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__23694\,
            I => \Inst_core.n1639\
        );

    \I__4593\ : InMux
    port map (
            O => \N__23687\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7913\
        );

    \I__4592\ : CascadeMux
    port map (
            O => \N__23684\,
            I => \N__23680\
        );

    \I__4591\ : InMux
    port map (
            O => \N__23683\,
            I => \N__23677\
        );

    \I__4590\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23674\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__23677\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__23674\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15\
        );

    \I__4587\ : CEMux
    port map (
            O => \N__23669\,
            I => \N__23665\
        );

    \I__4586\ : CEMux
    port map (
            O => \N__23668\,
            I => \N__23662\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__23665\,
            I => \N__23659\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__23662\,
            I => \N__23656\
        );

    \I__4583\ : Span4Mux_s3_v
    port map (
            O => \N__23659\,
            I => \N__23653\
        );

    \I__4582\ : Span4Mux_v
    port map (
            O => \N__23656\,
            I => \N__23650\
        );

    \I__4581\ : Span4Mux_s3_h
    port map (
            O => \N__23653\,
            I => \N__23647\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__23650\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4114\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__23647\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4114\
        );

    \I__4578\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23637\
        );

    \I__4577\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23634\
        );

    \I__4576\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23631\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__23637\,
            I => \N__23628\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__23634\,
            I => \N__23625\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__23631\,
            I => \Inst_core.configRegister_27\
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__23628\,
            I => \Inst_core.configRegister_27\
        );

    \I__4571\ : Odrv12
    port map (
            O => \N__23625\,
            I => \Inst_core.configRegister_27\
        );

    \I__4570\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23611\
        );

    \I__4568\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23608\
        );

    \I__4567\ : Odrv12
    port map (
            O => \N__23611\,
            I => \configRegister_7_adj_1353\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__23608\,
            I => \configRegister_7_adj_1353\
        );

    \I__4565\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23599\
        );

    \I__4564\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23596\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__23599\,
            I => \configRegister_11_adj_1349\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__23596\,
            I => \configRegister_11_adj_1349\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__23591\,
            I => \N__23588\
        );

    \I__4560\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23584\
        );

    \I__4559\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23581\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__23584\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__23581\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3\
        );

    \I__4556\ : InMux
    port map (
            O => \N__23576\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7901\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__4554\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23566\
        );

    \I__4553\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23563\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__23566\,
            I => \N__23560\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__23563\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4\
        );

    \I__4550\ : Odrv4
    port map (
            O => \N__23560\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4\
        );

    \I__4549\ : InMux
    port map (
            O => \N__23555\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7902\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__23552\,
            I => \N__23548\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__23551\,
            I => \N__23545\
        );

    \I__4546\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23542\
        );

    \I__4545\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23539\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__23542\,
            I => \N__23536\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__23539\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5\
        );

    \I__4542\ : Odrv4
    port map (
            O => \N__23536\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5\
        );

    \I__4541\ : InMux
    port map (
            O => \N__23531\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7903\
        );

    \I__4540\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23524\
        );

    \I__4539\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__23524\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__23521\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6\
        );

    \I__4536\ : InMux
    port map (
            O => \N__23516\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7904\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__23513\,
            I => \N__23509\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__23512\,
            I => \N__23506\
        );

    \I__4533\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23503\
        );

    \I__4532\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23500\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__23503\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__23500\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7\
        );

    \I__4529\ : InMux
    port map (
            O => \N__23495\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7905\
        );

    \I__4528\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23488\
        );

    \I__4527\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23485\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__23488\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__23485\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8\
        );

    \I__4524\ : InMux
    port map (
            O => \N__23480\,
            I => \bfn_8_3_0_\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__23477\,
            I => \N__23474\
        );

    \I__4522\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23470\
        );

    \I__4521\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23467\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__23470\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__23467\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9\
        );

    \I__4518\ : InMux
    port map (
            O => \N__23462\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7907\
        );

    \I__4517\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23455\
        );

    \I__4516\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23452\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__23455\,
            I => \configRegister_10_adj_1350\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23452\,
            I => \configRegister_10_adj_1350\
        );

    \I__4513\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23443\
        );

    \I__4512\ : InMux
    port map (
            O => \N__23446\,
            I => \N__23440\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__23443\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__23440\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10\
        );

    \I__4509\ : InMux
    port map (
            O => \N__23435\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7908\
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__4507\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23425\
        );

    \I__4506\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23422\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__23425\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__23422\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11\
        );

    \I__4503\ : InMux
    port map (
            O => \N__23417\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7909\
        );

    \I__4502\ : CascadeMux
    port map (
            O => \N__23414\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n8808_cascade_\
        );

    \I__4501\ : SRMux
    port map (
            O => \N__23411\,
            I => \N__23408\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__23408\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n3\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__23405\,
            I => \Inst_core.n1639_cascade_\
        );

    \I__4498\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__23399\,
            I => \Inst_core.n9054\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__4495\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23389\
        );

    \I__4494\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23386\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23389\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__23386\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0\
        );

    \I__4491\ : InMux
    port map (
            O => \N__23381\,
            I => \bfn_8_2_0_\
        );

    \I__4490\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__23375\,
            I => \N__23371\
        );

    \I__4488\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23368\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__23371\,
            I => \configRegister_1_adj_1359\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__23368\,
            I => \configRegister_1_adj_1359\
        );

    \I__4485\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23359\
        );

    \I__4484\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23356\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__23359\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__23356\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1\
        );

    \I__4481\ : InMux
    port map (
            O => \N__23351\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7899\
        );

    \I__4480\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23341\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23338\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__23341\,
            I => \configRegister_2_adj_1358\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__23338\,
            I => \configRegister_2_adj_1358\
        );

    \I__4475\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23329\
        );

    \I__4474\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23326\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__23329\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__23326\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2\
        );

    \I__4471\ : InMux
    port map (
            O => \N__23321\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7900\
        );

    \I__4470\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23311\
        );

    \I__4468\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23308\
        );

    \I__4467\ : Odrv12
    port map (
            O => \N__23311\,
            I => \configRegister_3_adj_1357\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__23308\,
            I => \configRegister_3_adj_1357\
        );

    \I__4465\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23299\
        );

    \I__4464\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23296\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__23299\,
            I => \N__23293\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__23296\,
            I => \N__23290\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__23293\,
            I => \N__23287\
        );

    \I__4460\ : Span12Mux_s11_h
    port map (
            O => \N__23290\,
            I => \N__23284\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__4458\ : Odrv12
    port map (
            O => \N__23284\,
            I => input_c_1
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__23281\,
            I => input_c_1
        );

    \I__4456\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23272\
        );

    \I__4455\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23269\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__23272\,
            I => \N__23266\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__23269\,
            I => \Inst_core.Inst_sync.synchronizedInput180_1\
        );

    \I__4452\ : Odrv4
    port map (
            O => \N__23266\,
            I => \Inst_core.Inst_sync.synchronizedInput180_1\
        );

    \I__4451\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__23258\,
            I => \N__23254\
        );

    \I__4449\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23251\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__23254\,
            I => \N__23246\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23246\
        );

    \I__4446\ : Span4Mux_h
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__23243\,
            I => input_c_2
        );

    \I__4444\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23234\
        );

    \I__4443\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23234\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__4441\ : Odrv4
    port map (
            O => \N__23231\,
            I => \Inst_core.Inst_sync.synchronizedInput180_2\
        );

    \I__4440\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23224\
        );

    \I__4439\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23221\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__23224\,
            I => \N__23218\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__23221\,
            I => \N__23215\
        );

    \I__4436\ : Span4Mux_h
    port map (
            O => \N__23218\,
            I => \N__23212\
        );

    \I__4435\ : Span4Mux_h
    port map (
            O => \N__23215\,
            I => \N__23209\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__23212\,
            I => input_c_3
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__23209\,
            I => input_c_3
        );

    \I__4432\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23200\
        );

    \I__4431\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23197\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__23200\,
            I => \N__23194\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__23197\,
            I => \Inst_core.Inst_sync.synchronizedInput180_3\
        );

    \I__4428\ : Odrv4
    port map (
            O => \N__23194\,
            I => \Inst_core.Inst_sync.synchronizedInput180_3\
        );

    \I__4427\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23185\
        );

    \I__4426\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23182\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23179\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__4423\ : IoSpan4Mux
    port map (
            O => \N__23179\,
            I => \N__23173\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__23176\,
            I => \N__23170\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__23173\,
            I => input_c_6
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__23170\,
            I => input_c_6
        );

    \I__4419\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23162\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__23162\,
            I => \N__23158\
        );

    \I__4417\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23155\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__23158\,
            I => \Inst_core.Inst_sync.synchronizedInput180_6\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__23155\,
            I => \Inst_core.Inst_sync.synchronizedInput180_6\
        );

    \I__4414\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23146\
        );

    \I__4413\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23143\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__23146\,
            I => \N__23140\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23137\
        );

    \I__4410\ : IoSpan4Mux
    port map (
            O => \N__23140\,
            I => \N__23134\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__23137\,
            I => \N__23131\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__23134\,
            I => input_c_5
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__23131\,
            I => input_c_5
        );

    \I__4406\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23123\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__23123\,
            I => \N__23119\
        );

    \I__4404\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23116\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__23119\,
            I => \Inst_core.Inst_sync.synchronizedInput180_5\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__23116\,
            I => \Inst_core.Inst_sync.synchronizedInput180_5\
        );

    \I__4401\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23107\
        );

    \I__4400\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23104\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__23107\,
            I => \Inst_core.Inst_sync.synchronizedInput180_7\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__23104\,
            I => \Inst_core.Inst_sync.synchronizedInput180_7\
        );

    \I__4397\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \Inst_core.n8518_cascade_\
        );

    \I__4396\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23093\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__23090\
        );

    \I__4394\ : Span12Mux_s10_v
    port map (
            O => \N__23090\,
            I => \N__23086\
        );

    \I__4393\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23083\
        );

    \I__4392\ : Odrv12
    port map (
            O => \N__23086\,
            I => \valueRegister_7_adj_1289\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__23083\,
            I => \valueRegister_7_adj_1289\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__23078\,
            I => \N__23075\
        );

    \I__4389\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__4387\ : Span4Mux_s2_v
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__4386\ : Span4Mux_h
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__4385\ : Span4Mux_v
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__23060\,
            I => \N__23057\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__23057\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_7\
        );

    \I__4382\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23050\
        );

    \I__4381\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23047\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__23050\,
            I => \N__23043\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__23047\,
            I => \N__23040\
        );

    \I__4378\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23033\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__23043\,
            I => \N__23030\
        );

    \I__4376\ : Span4Mux_h
    port map (
            O => \N__23040\,
            I => \N__23027\
        );

    \I__4375\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23022\
        );

    \I__4374\ : InMux
    port map (
            O => \N__23038\,
            I => \N__23019\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23015\
        );

    \I__4372\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23012\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__23033\,
            I => \N__23009\
        );

    \I__4370\ : Span4Mux_v
    port map (
            O => \N__23030\,
            I => \N__23006\
        );

    \I__4369\ : Sp12to4
    port map (
            O => \N__23027\,
            I => \N__23003\
        );

    \I__4368\ : InMux
    port map (
            O => \N__23026\,
            I => \N__23000\
        );

    \I__4367\ : InMux
    port map (
            O => \N__23025\,
            I => \N__22997\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__23022\,
            I => \N__22994\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__23019\,
            I => \N__22991\
        );

    \I__4364\ : InMux
    port map (
            O => \N__23018\,
            I => \N__22988\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__23015\,
            I => \N__22983\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__23012\,
            I => \N__22983\
        );

    \I__4361\ : Span4Mux_v
    port map (
            O => \N__23009\,
            I => \N__22980\
        );

    \I__4360\ : Span4Mux_v
    port map (
            O => \N__23006\,
            I => \N__22977\
        );

    \I__4359\ : Span12Mux_s5_v
    port map (
            O => \N__23003\,
            I => \N__22970\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22970\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22970\
        );

    \I__4356\ : Span4Mux_v
    port map (
            O => \N__22994\,
            I => \N__22965\
        );

    \I__4355\ : Span4Mux_h
    port map (
            O => \N__22991\,
            I => \N__22965\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__22988\,
            I => \memoryOut_7\
        );

    \I__4353\ : Odrv12
    port map (
            O => \N__22983\,
            I => \memoryOut_7\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__22980\,
            I => \memoryOut_7\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__22977\,
            I => \memoryOut_7\
        );

    \I__4350\ : Odrv12
    port map (
            O => \N__22970\,
            I => \memoryOut_7\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__22965\,
            I => \memoryOut_7\
        );

    \I__4348\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22948\
        );

    \I__4347\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22945\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__22948\,
            I => \N__22942\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__22945\,
            I => \N__22939\
        );

    \I__4344\ : Span4Mux_v
    port map (
            O => \N__22942\,
            I => \N__22936\
        );

    \I__4343\ : Odrv12
    port map (
            O => \N__22939\,
            I => \Inst_core.Inst_sync.demuxedInput_7\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__22936\,
            I => \Inst_core.Inst_sync.demuxedInput_7\
        );

    \I__4341\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22927\
        );

    \I__4340\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22924\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__22927\,
            I => \N__22921\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__22924\,
            I => \N__22917\
        );

    \I__4337\ : Span4Mux_v
    port map (
            O => \N__22921\,
            I => \N__22914\
        );

    \I__4336\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22911\
        );

    \I__4335\ : Span4Mux_h
    port map (
            O => \N__22917\,
            I => \N__22908\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__22914\,
            I => \N__22905\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22902\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__22908\,
            I => \Inst_core.Inst_sync.demuxedInput_2\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__22905\,
            I => \Inst_core.Inst_sync.demuxedInput_2\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__22902\,
            I => \Inst_core.Inst_sync.demuxedInput_2\
        );

    \I__4329\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22891\
        );

    \I__4328\ : InMux
    port map (
            O => \N__22894\,
            I => \N__22888\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__22891\,
            I => \N__22885\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__22888\,
            I => \N__22882\
        );

    \I__4325\ : Span4Mux_h
    port map (
            O => \N__22885\,
            I => \N__22879\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__22882\,
            I => \Inst_core.Inst_sync.demuxedInput_5\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__22879\,
            I => \Inst_core.Inst_sync.demuxedInput_5\
        );

    \I__4322\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22871\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__22868\,
            I => \Inst_core.Inst_sync.n9117\
        );

    \I__4319\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22861\
        );

    \I__4318\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22858\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__22861\,
            I => \N__22855\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__22858\,
            I => \N__22850\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__22855\,
            I => \N__22850\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__22850\,
            I => \N__22846\
        );

    \I__4313\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22843\
        );

    \I__4312\ : Span4Mux_v
    port map (
            O => \N__22846\,
            I => \N__22840\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__22843\,
            I => \N__22837\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__22840\,
            I => \Inst_core.Inst_sync.demuxedInput_3\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__22837\,
            I => \Inst_core.Inst_sync.demuxedInput_3\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__22832\,
            I => \N__22829\
        );

    \I__4307\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22824\
        );

    \I__4306\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22821\
        );

    \I__4305\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22818\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__22824\,
            I => \N__22815\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__22821\,
            I => \Inst_core.Inst_sync.synchronizedInput_5\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__22818\,
            I => \Inst_core.Inst_sync.synchronizedInput_5\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__22815\,
            I => \Inst_core.Inst_sync.synchronizedInput_5\
        );

    \I__4300\ : InMux
    port map (
            O => \N__22808\,
            I => \N__22796\
        );

    \I__4299\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22796\
        );

    \I__4298\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22791\
        );

    \I__4297\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22791\
        );

    \I__4296\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22788\
        );

    \I__4295\ : InMux
    port map (
            O => \N__22803\,
            I => \N__22785\
        );

    \I__4294\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22780\
        );

    \I__4293\ : InMux
    port map (
            O => \N__22801\,
            I => \N__22780\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__22796\,
            I => \N__22775\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22775\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__22788\,
            I => \Inst_core.Inst_sync.n2566\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__22785\,
            I => \Inst_core.Inst_sync.n2566\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__22780\,
            I => \Inst_core.Inst_sync.n2566\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__22775\,
            I => \Inst_core.Inst_sync.n2566\
        );

    \I__4286\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22754\
        );

    \I__4285\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22754\
        );

    \I__4284\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22754\
        );

    \I__4283\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22754\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__22754\,
            I => \N__22747\
        );

    \I__4281\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22742\
        );

    \I__4280\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22742\
        );

    \I__4279\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22739\
        );

    \I__4278\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22736\
        );

    \I__4277\ : Span4Mux_h
    port map (
            O => \N__22747\,
            I => \N__22733\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__22742\,
            I => \N__22730\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__22739\,
            I => \Inst_core.Inst_sync.n2564\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__22736\,
            I => \Inst_core.Inst_sync.n2564\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__22733\,
            I => \Inst_core.Inst_sync.n2564\
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__22730\,
            I => \Inst_core.Inst_sync.n2564\
        );

    \I__4271\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__4269\ : Odrv4
    port map (
            O => \N__22715\,
            I => \Inst_core.Inst_sync.n9129\
        );

    \I__4268\ : InMux
    port map (
            O => \N__22712\,
            I => \N__22708\
        );

    \I__4267\ : InMux
    port map (
            O => \N__22711\,
            I => \N__22704\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__22708\,
            I => \N__22701\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__22707\,
            I => \N__22698\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22693\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__22701\,
            I => \N__22693\
        );

    \I__4262\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22690\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__22693\,
            I => \Inst_core.Inst_sync.synchronizedInput_6\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__22690\,
            I => \Inst_core.Inst_sync.synchronizedInput_6\
        );

    \I__4259\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22682\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__22682\,
            I => \N__22678\
        );

    \I__4257\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22675\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__22678\,
            I => \N__22670\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__22675\,
            I => \N__22670\
        );

    \I__4254\ : Span4Mux_h
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__4253\ : IoSpan4Mux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__4252\ : Odrv4
    port map (
            O => \N__22664\,
            I => input_c_0
        );

    \I__4251\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22657\
        );

    \I__4250\ : InMux
    port map (
            O => \N__22660\,
            I => \N__22654\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__22657\,
            I => \N__22651\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__22654\,
            I => \Inst_core.Inst_sync.synchronizedInput180_0\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__22651\,
            I => \Inst_core.Inst_sync.synchronizedInput180_0\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__4245\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__4243\ : Span4Mux_h
    port map (
            O => \N__22637\,
            I => \N__22633\
        );

    \I__4242\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22630\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__22633\,
            I => \N__22627\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__22630\,
            I => \Inst_core.Inst_sync.filteredInput_0\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__22627\,
            I => \Inst_core.Inst_sync.filteredInput_0\
        );

    \I__4238\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22619\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__22619\,
            I => \Inst_core.Inst_sync.n2793\
        );

    \I__4236\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22612\
        );

    \I__4235\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22609\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__22612\,
            I => \N__22606\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__22609\,
            I => \flagInverted\
        );

    \I__4232\ : Odrv12
    port map (
            O => \N__22606\,
            I => \flagInverted\
        );

    \I__4231\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22589\
        );

    \I__4230\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22589\
        );

    \I__4229\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22589\
        );

    \I__4228\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22584\
        );

    \I__4227\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22584\
        );

    \I__4226\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22580\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__22589\,
            I => \N__22575\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__22584\,
            I => \N__22575\
        );

    \I__4223\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22572\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__22580\,
            I => \N__22569\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__22575\,
            I => \N__22566\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__22572\,
            I => \flagFilter\
        );

    \I__4219\ : Odrv12
    port map (
            O => \N__22569\,
            I => \flagFilter\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__22566\,
            I => \flagFilter\
        );

    \I__4217\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22555\
        );

    \I__4216\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22552\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__22555\,
            I => \N__22549\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__22552\,
            I => \N__22543\
        );

    \I__4213\ : Span4Mux_h
    port map (
            O => \N__22549\,
            I => \N__22543\
        );

    \I__4212\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22540\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__22543\,
            I => \Inst_core.Inst_sync.demuxedInput_1\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__22540\,
            I => \Inst_core.Inst_sync.demuxedInput_1\
        );

    \I__4209\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__22532\,
            I => \Inst_core.Inst_sync.n2787\
        );

    \I__4207\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__22526\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_5\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__22523\,
            I => \N__22520\
        );

    \I__4204\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22517\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__22517\,
            I => \syncedInput_6\
        );

    \I__4202\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__22505\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_6\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__4197\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__22496\,
            I => \syncedInput_3\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__4194\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22487\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__4192\ : Span4Mux_h
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__22481\,
            I => \syncedInput_7\
        );

    \I__4190\ : InMux
    port map (
            O => \N__22478\,
            I => \N__22474\
        );

    \I__4189\ : InMux
    port map (
            O => \N__22477\,
            I => \N__22471\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__22474\,
            I => \valueRegister_7_adj_1329\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__22471\,
            I => \valueRegister_7_adj_1329\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__22466\,
            I => \N__22463\
        );

    \I__4185\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22457\
        );

    \I__4183\ : Span4Mux_v
    port map (
            O => \N__22457\,
            I => \N__22453\
        );

    \I__4182\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22450\
        );

    \I__4181\ : Span4Mux_h
    port map (
            O => \N__22453\,
            I => \N__22447\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__22450\,
            I => \Inst_core.Inst_sync.filteredInput_1\
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__22447\,
            I => \Inst_core.Inst_sync.filteredInput_1\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__4177\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__22436\,
            I => \N__22432\
        );

    \I__4175\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22429\
        );

    \I__4174\ : Span12Mux_s7_h
    port map (
            O => \N__22432\,
            I => \N__22426\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__22429\,
            I => \Inst_core.Inst_sync.filteredInput_3\
        );

    \I__4172\ : Odrv12
    port map (
            O => \N__22426\,
            I => \Inst_core.Inst_sync.filteredInput_3\
        );

    \I__4171\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__22418\,
            I => \Inst_core.Inst_sync.n2791\
        );

    \I__4169\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__4167\ : Span4Mux_s2_h
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__22403\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_1\
        );

    \I__4164\ : SRMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__4162\ : Span4Mux_v
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__22391\,
            I => \N__22388\
        );

    \I__4160\ : Span4Mux_h
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__22385\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4746\
        );

    \I__4158\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__22379\,
            I => \N__22375\
        );

    \I__4156\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22372\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__22375\,
            I => \N__22369\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__22372\,
            I => fwd_15
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__22369\,
            I => fwd_15
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__22364\,
            I => \Inst_core.Inst_controller.n22_cascade_\
        );

    \I__4151\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22357\
        );

    \I__4150\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22354\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__22357\,
            I => fwd_6
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__22354\,
            I => fwd_6
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__22349\,
            I => \Inst_core.Inst_controller.n4_adj_986_cascade_\
        );

    \I__4146\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22342\
        );

    \I__4145\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22339\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__22342\,
            I => fwd_5
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__22339\,
            I => fwd_5
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__22334\,
            I => \Inst_core.Inst_controller.n4_adj_987_cascade_\
        );

    \I__4141\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__22328\,
            I => \Inst_core.Inst_controller.n8486\
        );

    \I__4139\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__4137\ : Span4Mux_h
    port map (
            O => \N__22319\,
            I => \N__22314\
        );

    \I__4136\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22311\
        );

    \I__4135\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22308\
        );

    \I__4134\ : Span4Mux_v
    port map (
            O => \N__22314\,
            I => \N__22305\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22302\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__22308\,
            I => \Inst_core.Inst_sync.demuxedInput_0\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__22305\,
            I => \Inst_core.Inst_sync.demuxedInput_0\
        );

    \I__4130\ : Odrv12
    port map (
            O => \N__22302\,
            I => \Inst_core.Inst_sync.demuxedInput_0\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22286\
        );

    \I__4127\ : InMux
    port map (
            O => \N__22291\,
            I => \N__22286\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__22286\,
            I => \N__22282\
        );

    \I__4125\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22279\
        );

    \I__4124\ : Span4Mux_s3_h
    port map (
            O => \N__22282\,
            I => \N__22272\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22272\
        );

    \I__4122\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22269\
        );

    \I__4121\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22266\
        );

    \I__4120\ : Span4Mux_h
    port map (
            O => \N__22272\,
            I => \N__22261\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__22269\,
            I => \N__22261\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__22266\,
            I => \N__22257\
        );

    \I__4117\ : Span4Mux_v
    port map (
            O => \N__22261\,
            I => \N__22253\
        );

    \I__4116\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22250\
        );

    \I__4115\ : Sp12to4
    port map (
            O => \N__22257\,
            I => \N__22247\
        );

    \I__4114\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22244\
        );

    \I__4113\ : Sp12to4
    port map (
            O => \N__22253\,
            I => \N__22239\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22239\
        );

    \I__4111\ : Span12Mux_s11_v
    port map (
            O => \N__22247\,
            I => \N__22236\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__22244\,
            I => \N__22231\
        );

    \I__4109\ : Span12Mux_s8_h
    port map (
            O => \N__22239\,
            I => \N__22231\
        );

    \I__4108\ : Odrv12
    port map (
            O => \N__22236\,
            I => \wrFlags\
        );

    \I__4107\ : Odrv12
    port map (
            O => \N__22231\,
            I => \wrFlags\
        );

    \I__4106\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22220\
        );

    \I__4105\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22220\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__22220\,
            I => \N__22213\
        );

    \I__4103\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22210\
        );

    \I__4102\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22207\
        );

    \I__4101\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22204\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__22216\,
            I => \N__22200\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__22213\,
            I => \N__22197\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__22210\,
            I => \N__22194\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__22207\,
            I => \N__22189\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__22204\,
            I => \N__22189\
        );

    \I__4095\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22186\
        );

    \I__4094\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22183\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__22197\,
            I => cmd_32
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__22194\,
            I => cmd_32
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__22189\,
            I => cmd_32
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__22186\,
            I => cmd_32
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__22183\,
            I => cmd_32
        );

    \I__4088\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22168\
        );

    \I__4087\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22165\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22162\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__22165\,
            I => \N__22158\
        );

    \I__4084\ : Span4Mux_s2_h
    port map (
            O => \N__22162\,
            I => \N__22155\
        );

    \I__4083\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22152\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__22158\,
            I => \N__22147\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__22155\,
            I => \N__22147\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__22152\,
            I => \configRegister_20\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__22147\,
            I => \configRegister_20\
        );

    \I__4078\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__22136\,
            I => \N__22132\
        );

    \I__4075\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22129\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__22132\,
            I => \valueRegister_1_adj_1295\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__22129\,
            I => \valueRegister_1_adj_1295\
        );

    \I__4072\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22119\
        );

    \I__4071\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22114\
        );

    \I__4070\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22114\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__22119\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__22114\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1\
        );

    \I__4067\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22103\
        );

    \I__4066\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22103\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__22103\,
            I => \N__22099\
        );

    \I__4064\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22096\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__22099\,
            I => \N__22093\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__22096\,
            I => \configRegister_22_adj_1340\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__22093\,
            I => \configRegister_22_adj_1340\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__22088\,
            I => \N__22083\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__22087\,
            I => \N__22080\
        );

    \I__4058\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22075\
        );

    \I__4057\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22075\
        );

    \I__4056\ : InMux
    port map (
            O => \N__22080\,
            I => \N__22071\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__22075\,
            I => \N__22068\
        );

    \I__4054\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22065\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__22071\,
            I => \N__22062\
        );

    \I__4052\ : Span4Mux_v
    port map (
            O => \N__22068\,
            I => \N__22058\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__22065\,
            I => \N__22053\
        );

    \I__4050\ : Span4Mux_v
    port map (
            O => \N__22062\,
            I => \N__22053\
        );

    \I__4049\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22050\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__22058\,
            I => \N__22047\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__22053\,
            I => \N__22044\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__22050\,
            I => \configRegister_21\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__22047\,
            I => \configRegister_21\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__22044\,
            I => \configRegister_21\
        );

    \I__4043\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22031\
        );

    \I__4042\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22028\
        );

    \I__4041\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22019\
        );

    \I__4040\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22019\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__22031\,
            I => \N__22016\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22013\
        );

    \I__4037\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22010\
        );

    \I__4036\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22007\
        );

    \I__4035\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22004\
        );

    \I__4034\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22001\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__21998\
        );

    \I__4032\ : Span4Mux_h
    port map (
            O => \N__22016\,
            I => \N__21995\
        );

    \I__4031\ : Span4Mux_h
    port map (
            O => \N__22013\,
            I => \N__21992\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__21985\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__22007\,
            I => \N__21985\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__22004\,
            I => \N__21985\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21982\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__21998\,
            I => \N__21979\
        );

    \I__4025\ : Span4Mux_s3_h
    port map (
            O => \N__21995\,
            I => \N__21976\
        );

    \I__4024\ : Span4Mux_v
    port map (
            O => \N__21992\,
            I => \N__21971\
        );

    \I__4023\ : Span4Mux_v
    port map (
            O => \N__21985\,
            I => \N__21971\
        );

    \I__4022\ : Span12Mux_s8_h
    port map (
            O => \N__21982\,
            I => \N__21964\
        );

    \I__4021\ : Sp12to4
    port map (
            O => \N__21979\,
            I => \N__21964\
        );

    \I__4020\ : Sp12to4
    port map (
            O => \N__21976\,
            I => \N__21964\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__21971\,
            I => wrtrigmask_1
        );

    \I__4018\ : Odrv12
    port map (
            O => \N__21964\,
            I => wrtrigmask_1
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__21959\,
            I => \N__21953\
        );

    \I__4016\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21943\
        );

    \I__4015\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21943\
        );

    \I__4014\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21943\
        );

    \I__4013\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21943\
        );

    \I__4012\ : InMux
    port map (
            O => \N__21952\,
            I => \N__21940\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__21943\,
            I => \N__21937\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__21940\,
            I => \configRegister_21_adj_1341\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__21937\,
            I => \configRegister_21_adj_1341\
        );

    \I__4008\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21926\
        );

    \I__4007\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21926\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__21926\,
            I => \N__21922\
        );

    \I__4005\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21919\
        );

    \I__4004\ : Span4Mux_v
    port map (
            O => \N__21922\,
            I => \N__21916\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__21919\,
            I => \configRegister_22_adj_1380\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__21916\,
            I => \configRegister_22_adj_1380\
        );

    \I__4001\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21905\
        );

    \I__4000\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21905\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21901\
        );

    \I__3998\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21898\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__21901\,
            I => \N__21895\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__21898\,
            I => \configRegister_23\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__21895\,
            I => \configRegister_23\
        );

    \I__3994\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21881\
        );

    \I__3993\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21878\
        );

    \I__3992\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21875\
        );

    \I__3991\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21866\
        );

    \I__3990\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21866\
        );

    \I__3989\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21866\
        );

    \I__3988\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21866\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21862\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__21878\,
            I => \N__21859\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21856\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21853\
        );

    \I__3983\ : InMux
    port map (
            O => \N__21865\,
            I => \N__21850\
        );

    \I__3982\ : Span4Mux_h
    port map (
            O => \N__21862\,
            I => \N__21847\
        );

    \I__3981\ : Span4Mux_s3_h
    port map (
            O => \N__21859\,
            I => \N__21842\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__21856\,
            I => \N__21842\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__21853\,
            I => \N__21837\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21837\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__21847\,
            I => wrtrigmask_0
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__21842\,
            I => wrtrigmask_0
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__21837\,
            I => wrtrigmask_0
        );

    \I__3974\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21826\
        );

    \I__3973\ : InMux
    port map (
            O => \N__21829\,
            I => \N__21823\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__21826\,
            I => \maskRegister_0\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__21823\,
            I => \maskRegister_0\
        );

    \I__3970\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21811\
        );

    \I__3969\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21811\
        );

    \I__3968\ : InMux
    port map (
            O => \N__21816\,
            I => \N__21808\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21805\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__21808\,
            I => \configRegister_20_adj_1382\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__21805\,
            I => \configRegister_20_adj_1382\
        );

    \I__3964\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__21797\,
            I => \N__21793\
        );

    \I__3962\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21790\
        );

    \I__3961\ : Odrv12
    port map (
            O => \N__21793\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__21790\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6\
        );

    \I__3959\ : CascadeMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__3958\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__21776\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_7\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__3954\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__21767\,
            I => \N__21763\
        );

    \I__3952\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21760\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__21763\,
            I => \configRegister_15_adj_1385\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__21760\,
            I => \configRegister_15_adj_1385\
        );

    \I__3949\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21751\
        );

    \I__3948\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21748\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__21751\,
            I => \configRegister_24_adj_1378\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__21748\,
            I => \configRegister_24_adj_1378\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__21743\,
            I => \N__21738\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__21742\,
            I => \N__21735\
        );

    \I__3943\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21716\
        );

    \I__3942\ : InMux
    port map (
            O => \N__21738\,
            I => \N__21716\
        );

    \I__3941\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21716\
        );

    \I__3940\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21716\
        );

    \I__3939\ : InMux
    port map (
            O => \N__21733\,
            I => \N__21716\
        );

    \I__3938\ : InMux
    port map (
            O => \N__21732\,
            I => \N__21716\
        );

    \I__3937\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21713\
        );

    \I__3936\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21708\
        );

    \I__3935\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21708\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21705\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__21713\,
            I => \N__21702\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__21708\,
            I => \N__21699\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__21705\,
            I => \N__21694\
        );

    \I__3930\ : Span4Mux_h
    port map (
            O => \N__21702\,
            I => \N__21694\
        );

    \I__3929\ : Span4Mux_s3_h
    port map (
            O => \N__21699\,
            I => \N__21691\
        );

    \I__3928\ : Span4Mux_v
    port map (
            O => \N__21694\,
            I => \N__21688\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__21691\,
            I => \Inst_eia232.Inst_transmitter.n4246\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__21688\,
            I => \Inst_eia232.Inst_transmitter.n4246\
        );

    \I__3925\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21678\
        );

    \I__3924\ : CEMux
    port map (
            O => \N__21682\,
            I => \N__21673\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21670\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__21678\,
            I => \N__21659\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__21677\,
            I => \N__21652\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__21676\,
            I => \N__21649\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__21673\,
            I => \N__21646\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21643\
        );

    \I__3917\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21638\
        );

    \I__3916\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21638\
        );

    \I__3915\ : InMux
    port map (
            O => \N__21667\,
            I => \N__21633\
        );

    \I__3914\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21633\
        );

    \I__3913\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21624\
        );

    \I__3912\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21624\
        );

    \I__3911\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21624\
        );

    \I__3910\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21624\
        );

    \I__3909\ : Span4Mux_h
    port map (
            O => \N__21659\,
            I => \N__21621\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__21658\,
            I => \N__21618\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__21657\,
            I => \N__21615\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__21656\,
            I => \N__21612\
        );

    \I__3905\ : CEMux
    port map (
            O => \N__21655\,
            I => \N__21607\
        );

    \I__3904\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21602\
        );

    \I__3903\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21602\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__21646\,
            I => \N__21599\
        );

    \I__3901\ : Span4Mux_h
    port map (
            O => \N__21643\,
            I => \N__21596\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__21638\,
            I => \N__21587\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__21633\,
            I => \N__21587\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__21624\,
            I => \N__21587\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__21621\,
            I => \N__21587\
        );

    \I__3896\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21584\
        );

    \I__3895\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21575\
        );

    \I__3894\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21575\
        );

    \I__3893\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21575\
        );

    \I__3892\ : InMux
    port map (
            O => \N__21610\,
            I => \N__21575\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__21607\,
            I => \N__21570\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__21602\,
            I => \N__21570\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__21599\,
            I => \N__21565\
        );

    \I__3888\ : Span4Mux_v
    port map (
            O => \N__21596\,
            I => \N__21565\
        );

    \I__3887\ : Span4Mux_v
    port map (
            O => \N__21587\,
            I => \N__21562\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__21584\,
            I => n4005
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__21575\,
            I => n4005
        );

    \I__3884\ : Odrv12
    port map (
            O => \N__21570\,
            I => n4005
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__21565\,
            I => n4005
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__21562\,
            I => n4005
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__3880\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21542\
        );

    \I__3879\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21542\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__21542\,
            I => \disabledGroupsReg_0\
        );

    \I__3877\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21536\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__3875\ : Span4Mux_s2_h
    port map (
            O => \N__21533\,
            I => \N__21529\
        );

    \I__3874\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21526\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__21529\,
            I => \N__21523\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__21526\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_0\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__21523\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_0\
        );

    \I__3870\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21514\
        );

    \I__3869\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21511\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__21514\,
            I => \configRegister_11_adj_1389\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__21511\,
            I => \configRegister_11_adj_1389\
        );

    \I__3866\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21502\
        );

    \I__3865\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21499\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__21502\,
            I => \configRegister_10_adj_1390\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__21499\,
            I => \configRegister_10_adj_1390\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__3861\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__21488\,
            I => \N__21484\
        );

    \I__3859\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21481\
        );

    \I__3858\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21478\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__21481\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__21478\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16\
        );

    \I__3855\ : InMux
    port map (
            O => \N__21473\,
            I => \N__21467\
        );

    \I__3854\ : InMux
    port map (
            O => \N__21472\,
            I => \N__21467\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__21467\,
            I => \N__21463\
        );

    \I__3852\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21460\
        );

    \I__3851\ : Span4Mux_h
    port map (
            O => \N__21463\,
            I => \N__21457\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__21460\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__21457\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__21452\,
            I => \N__21449\
        );

    \I__3847\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21445\
        );

    \I__3846\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21442\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__21445\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__21442\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6\
        );

    \I__3843\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21433\
        );

    \I__3842\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21430\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__21433\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__21430\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1\
        );

    \I__3839\ : CascadeMux
    port map (
            O => \N__21425\,
            I => \N__21421\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__21424\,
            I => \N__21418\
        );

    \I__3837\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21415\
        );

    \I__3836\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21412\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__21415\,
            I => \N__21409\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__21412\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__21409\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__3831\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21397\
        );

    \I__3830\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21394\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__21397\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__21394\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0\
        );

    \I__3827\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21386\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__21386\,
            I => \N__21383\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__21380\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n28\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__21377\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n25_cascade_\
        );

    \I__3822\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__3820\ : Span4Mux_h
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__21365\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n27\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__3817\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21355\
        );

    \I__3816\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21352\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__21355\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__21352\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13\
        );

    \I__3813\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21343\
        );

    \I__3812\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21340\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__21343\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__21340\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__21335\,
            I => \N__21331\
        );

    \I__3808\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21328\
        );

    \I__3807\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21325\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__21328\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__21325\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5\
        );

    \I__3804\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21316\
        );

    \I__3803\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21313\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__21316\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__21313\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8\
        );

    \I__3800\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__21305\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n26\
        );

    \I__3798\ : InMux
    port map (
            O => \N__21302\,
            I => \N__21299\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__21299\,
            I => \N__21295\
        );

    \I__3796\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21292\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__21295\,
            I => \valueRegister_6_adj_1370\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__21292\,
            I => \valueRegister_6_adj_1370\
        );

    \I__3793\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21283\
        );

    \I__3792\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21280\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__21283\,
            I => \configRegister_5_adj_1395\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__21280\,
            I => \configRegister_5_adj_1395\
        );

    \I__3789\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21271\
        );

    \I__3788\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21268\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__21271\,
            I => \valueRegister_7_adj_1369\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__21268\,
            I => \valueRegister_7_adj_1369\
        );

    \I__3785\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__21260\,
            I => \N__21256\
        );

    \I__3783\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21253\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__21256\,
            I => \N__21248\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__21253\,
            I => \N__21248\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__21245\,
            I => input_c_4
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__21242\,
            I => \N__21238\
        );

    \I__3777\ : InMux
    port map (
            O => \N__21241\,
            I => \N__21235\
        );

    \I__3776\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21232\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__21235\,
            I => \Inst_core.Inst_sync.synchronizedInput180_4\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__21232\,
            I => \Inst_core.Inst_sync.synchronizedInput180_4\
        );

    \I__3773\ : SRMux
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__3771\ : Span4Mux_s2_v
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__21218\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4765\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__21215\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n25_cascade_\
        );

    \I__3768\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__21209\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n27\
        );

    \I__3766\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__21203\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n26\
        );

    \I__3764\ : SRMux
    port map (
            O => \N__21200\,
            I => \N__21197\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__3762\ : Span4Mux_v
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__3761\ : Span4Mux_h
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__21188\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4766\
        );

    \I__3759\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__21182\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n28\
        );

    \I__3757\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21175\
        );

    \I__3756\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21172\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__21175\,
            I => \N__21169\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__21172\,
            I => \Inst_core.Inst_sync.filteredInput_5\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__21169\,
            I => \Inst_core.Inst_sync.filteredInput_5\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__21164\,
            I => \Inst_core.Inst_sync.n9063_cascade_\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__3750\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21155\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__21155\,
            I => \syncedInput_5\
        );

    \I__3748\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21148\
        );

    \I__3747\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21145\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__21148\,
            I => \N__21139\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__21145\,
            I => \N__21139\
        );

    \I__3744\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21136\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__21139\,
            I => \Inst_core.Inst_sync.synchronizedInput_4\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__21136\,
            I => \Inst_core.Inst_sync.synchronizedInput_4\
        );

    \I__3741\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21128\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__3739\ : Span4Mux_h
    port map (
            O => \N__21125\,
            I => \N__21121\
        );

    \I__3738\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21118\
        );

    \I__3737\ : Span4Mux_s1_v
    port map (
            O => \N__21121\,
            I => \N__21115\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__21118\,
            I => \Inst_core.Inst_sync.filteredInput_4\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__21115\,
            I => \Inst_core.Inst_sync.filteredInput_4\
        );

    \I__3734\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21106\
        );

    \I__3733\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21103\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__21106\,
            I => \Inst_core.Inst_sync.demuxedInput_4\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__21103\,
            I => \Inst_core.Inst_sync.demuxedInput_4\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__21098\,
            I => \Inst_core.Inst_sync.n9057_cascade_\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__3728\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__21089\,
            I => \syncedInput_4\
        );

    \I__3726\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__21083\,
            I => \Inst_core.Inst_sync.Inst_filter.input180Delay_6\
        );

    \I__3724\ : SRMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__3722\ : Span4Mux_h
    port map (
            O => \N__21074\,
            I => \N__21071\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__21071\,
            I => \N__21068\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__21068\,
            I => \Inst_core.Inst_sync.Inst_filter.n4734\
        );

    \I__3719\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21062\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__21062\,
            I => \Inst_core.Inst_sync.Inst_filter.input180Delay_5\
        );

    \I__3717\ : SRMux
    port map (
            O => \N__21059\,
            I => \N__21056\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__21056\,
            I => \N__21053\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__21050\,
            I => \Inst_core.Inst_sync.Inst_filter.n4733\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__3712\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__21041\,
            I => \N__21037\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21034\
        );

    \I__3709\ : Span4Mux_v
    port map (
            O => \N__21037\,
            I => \N__21031\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__21034\,
            I => \Inst_core.Inst_sync.filteredInput_2\
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__21031\,
            I => \Inst_core.Inst_sync.filteredInput_2\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__21026\,
            I => \Inst_core.Inst_sync.n2789_cascade_\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__21023\,
            I => \N__21020\
        );

    \I__3704\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__21017\,
            I => \syncedInput_2\
        );

    \I__3702\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__21007\
        );

    \I__3700\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21004\
        );

    \I__3699\ : Span4Mux_v
    port map (
            O => \N__21007\,
            I => \N__21001\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__21004\,
            I => \Inst_core.Inst_sync.demuxedInput_6\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__21001\,
            I => \Inst_core.Inst_sync.demuxedInput_6\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__20996\,
            I => \N__20992\
        );

    \I__3695\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20989\
        );

    \I__3694\ : InMux
    port map (
            O => \N__20992\,
            I => \N__20986\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__20989\,
            I => \Inst_core.Inst_sync.filteredInput_6\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__20986\,
            I => \Inst_core.Inst_sync.filteredInput_6\
        );

    \I__3691\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20977\
        );

    \I__3690\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20974\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__20977\,
            I => \maskRegister_4_adj_1284\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__20974\,
            I => \maskRegister_4_adj_1284\
        );

    \I__3687\ : SRMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__20966\,
            I => \N__20963\
        );

    \I__3685\ : Sp12to4
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__3684\ : Odrv12
    port map (
            O => \N__20960\,
            I => \Inst_core.Inst_sync.Inst_filter.n4637\
        );

    \I__3683\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20953\
        );

    \I__3682\ : InMux
    port map (
            O => \N__20956\,
            I => \N__20950\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20947\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__20950\,
            I => \maskRegister_1\
        );

    \I__3679\ : Odrv12
    port map (
            O => \N__20947\,
            I => \maskRegister_1\
        );

    \I__3678\ : SRMux
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__3676\ : Span4Mux_v
    port map (
            O => \N__20936\,
            I => \N__20933\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__20933\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4739\
        );

    \I__3674\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__20927\,
            I => \Inst_core.Inst_sync.Inst_filter.input180Delay_7\
        );

    \I__3672\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20920\
        );

    \I__3671\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20917\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20914\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__20917\,
            I => \maskRegister_1_adj_1287\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__20914\,
            I => \maskRegister_1_adj_1287\
        );

    \I__3667\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20905\
        );

    \I__3666\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20902\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__20905\,
            I => \maskRegister_2_adj_1286\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__20902\,
            I => \maskRegister_2_adj_1286\
        );

    \I__3663\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20893\
        );

    \I__3662\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__20893\,
            I => \N__20887\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__20890\,
            I => \maskRegister_3_adj_1285\
        );

    \I__3659\ : Odrv12
    port map (
            O => \N__20887\,
            I => \maskRegister_3_adj_1285\
        );

    \I__3658\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20875\
        );

    \I__3656\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20872\
        );

    \I__3655\ : Span4Mux_v
    port map (
            O => \N__20875\,
            I => \N__20869\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__20872\,
            I => \maskRegister_5_adj_1283\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__20869\,
            I => \maskRegister_5_adj_1283\
        );

    \I__3652\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20859\
        );

    \I__3651\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20854\
        );

    \I__3650\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20854\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__20859\,
            I => \configRegister_20_adj_1302\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__20854\,
            I => \configRegister_20_adj_1302\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__3646\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20842\
        );

    \I__3645\ : InMux
    port map (
            O => \N__20845\,
            I => \N__20839\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__20842\,
            I => \configRegister_24_adj_1298\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__20839\,
            I => \configRegister_24_adj_1298\
        );

    \I__3642\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20830\
        );

    \I__3641\ : InMux
    port map (
            O => \N__20833\,
            I => \N__20827\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__20830\,
            I => \N__20824\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__20827\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__20824\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__20819\,
            I => \N__20814\
        );

    \I__3636\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20809\
        );

    \I__3635\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20809\
        );

    \I__3634\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20806\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__20809\,
            I => \N__20803\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__20806\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__20803\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16\
        );

    \I__3630\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20794\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__20797\,
            I => \N__20791\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__20794\,
            I => \N__20787\
        );

    \I__3627\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20782\
        );

    \I__3626\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20782\
        );

    \I__3625\ : Odrv12
    port map (
            O => \N__20787\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__20782\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__20777\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_cascade_\
        );

    \I__3622\ : InMux
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__20771\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9078\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__20768\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_cascade_\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__20765\,
            I => \N__20758\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__20764\,
            I => \N__20755\
        );

    \I__3617\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20752\
        );

    \I__3616\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20743\
        );

    \I__3615\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20743\
        );

    \I__3614\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20743\
        );

    \I__3613\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20743\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__20752\,
            I => \configRegister_21_adj_1301\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__20743\,
            I => \configRegister_21_adj_1301\
        );

    \I__3610\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20733\
        );

    \I__3609\ : InMux
    port map (
            O => \N__20737\,
            I => \N__20728\
        );

    \I__3608\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20728\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__20733\,
            I => \configRegister_23_adj_1299\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__20728\,
            I => \configRegister_23_adj_1299\
        );

    \I__3605\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20716\
        );

    \I__3604\ : InMux
    port map (
            O => \N__20722\,
            I => \N__20716\
        );

    \I__3603\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20713\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20710\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__20713\,
            I => \configRegister_22_adj_1300\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__20710\,
            I => \configRegister_22_adj_1300\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__20705\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9072_cascade_\
        );

    \I__3598\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20696\
        );

    \I__3597\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20692\
        );

    \I__3596\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20684\
        );

    \I__3595\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20684\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__20696\,
            I => \N__20681\
        );

    \I__3593\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20678\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__20692\,
            I => \N__20675\
        );

    \I__3591\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20672\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__20690\,
            I => \N__20669\
        );

    \I__3589\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20666\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__20684\,
            I => \N__20663\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__20681\,
            I => \N__20654\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__20678\,
            I => \N__20654\
        );

    \I__3585\ : Span4Mux_s3_v
    port map (
            O => \N__20675\,
            I => \N__20654\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__20672\,
            I => \N__20654\
        );

    \I__3583\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20651\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20644\
        );

    \I__3581\ : Span4Mux_v
    port map (
            O => \N__20663\,
            I => \N__20644\
        );

    \I__3580\ : Span4Mux_v
    port map (
            O => \N__20654\,
            I => \N__20644\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__20651\,
            I => \N__20641\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__20644\,
            I => \N__20638\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__20641\,
            I => wrtrigval_0
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__20638\,
            I => wrtrigval_0
        );

    \I__3575\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__20630\,
            I => \N__20625\
        );

    \I__3573\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20620\
        );

    \I__3572\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20620\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__20625\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__20620\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1\
        );

    \I__3569\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20611\
        );

    \I__3568\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20608\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__20611\,
            I => \valueRegister_1\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__20608\,
            I => \valueRegister_1\
        );

    \I__3565\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20599\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__20602\,
            I => \N__20594\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__20599\,
            I => \N__20590\
        );

    \I__3562\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20587\
        );

    \I__3561\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20584\
        );

    \I__3560\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20581\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__20593\,
            I => \N__20577\
        );

    \I__3558\ : Span4Mux_s2_v
    port map (
            O => \N__20590\,
            I => \N__20571\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__20587\,
            I => \N__20571\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__20584\,
            I => \N__20568\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20565\
        );

    \I__3554\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20562\
        );

    \I__3553\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20558\
        );

    \I__3552\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20555\
        );

    \I__3551\ : Span4Mux_v
    port map (
            O => \N__20571\,
            I => \N__20551\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__20568\,
            I => \N__20546\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__20565\,
            I => \N__20546\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__20562\,
            I => \N__20543\
        );

    \I__3547\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20540\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__20558\,
            I => \N__20535\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20535\
        );

    \I__3544\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20532\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__20551\,
            I => \configRegister_26\
        );

    \I__3542\ : Odrv4
    port map (
            O => \N__20546\,
            I => \configRegister_26\
        );

    \I__3541\ : Odrv12
    port map (
            O => \N__20543\,
            I => \configRegister_26\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__20540\,
            I => \configRegister_26\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__20535\,
            I => \configRegister_26\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__20532\,
            I => \configRegister_26\
        );

    \I__3537\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20516\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__3535\ : Span4Mux_v
    port map (
            O => \N__20513\,
            I => \N__20510\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__20510\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_1\
        );

    \I__3533\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20504\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20501\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__20501\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_3\
        );

    \I__3530\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20494\
        );

    \I__3529\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20491\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__20494\,
            I => \N__20488\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__20491\,
            I => \configRegister_0_adj_1400\
        );

    \I__3526\ : Odrv12
    port map (
            O => \N__20488\,
            I => \configRegister_0_adj_1400\
        );

    \I__3525\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20476\
        );

    \I__3524\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20476\
        );

    \I__3523\ : InMux
    port map (
            O => \N__20481\,
            I => \N__20473\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__20476\,
            I => \N__20470\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__20473\,
            I => \configRegister_20_adj_1342\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__20470\,
            I => \configRegister_20_adj_1342\
        );

    \I__3519\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20458\
        );

    \I__3517\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20455\
        );

    \I__3516\ : Span4Mux_s3_v
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__20455\,
            I => \configRegister_4_adj_1396\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__20452\,
            I => \configRegister_4_adj_1396\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__20447\,
            I => \N__20442\
        );

    \I__3512\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20439\
        );

    \I__3511\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20436\
        );

    \I__3510\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20433\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__20439\,
            I => \N__20428\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20428\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__20433\,
            I => cmd_39
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__20428\,
            I => cmd_39
        );

    \I__3505\ : SRMux
    port map (
            O => \N__20423\,
            I => \N__20420\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__3503\ : Odrv12
    port map (
            O => \N__20417\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4641\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__20414\,
            I => \N__20407\
        );

    \I__3501\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20404\
        );

    \I__3500\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20395\
        );

    \I__3499\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20395\
        );

    \I__3498\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20395\
        );

    \I__3497\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20395\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__20404\,
            I => \configRegister_21_adj_1381\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__20395\,
            I => \configRegister_21_adj_1381\
        );

    \I__3494\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20386\
        );

    \I__3493\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20383\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__20386\,
            I => \maskRegister_6_adj_1362\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__20383\,
            I => \maskRegister_6_adj_1362\
        );

    \I__3490\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20374\
        );

    \I__3489\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20371\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__20374\,
            I => \maskRegister_7_adj_1361\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__20371\,
            I => \maskRegister_7_adj_1361\
        );

    \I__3486\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20362\
        );

    \I__3485\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20359\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__20362\,
            I => \maskRegister_4_adj_1364\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__20359\,
            I => \maskRegister_4_adj_1364\
        );

    \I__3482\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__3480\ : Span4Mux_s2_v
    port map (
            O => \N__20348\,
            I => \N__20344\
        );

    \I__3479\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20341\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__20344\,
            I => \configRegister_6_adj_1394\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__20341\,
            I => \configRegister_6_adj_1394\
        );

    \I__3476\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20332\
        );

    \I__3475\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20329\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__20332\,
            I => \maskRegister_3_adj_1365\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__20329\,
            I => \maskRegister_3_adj_1365\
        );

    \I__3472\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__20321\,
            I => \N__20317\
        );

    \I__3470\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20314\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__20317\,
            I => \configRegister_7_adj_1393\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__20314\,
            I => \configRegister_7_adj_1393\
        );

    \I__3467\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20306\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__3465\ : Span4Mux_s3_h
    port map (
            O => \N__20303\,
            I => \N__20300\
        );

    \I__3464\ : Span4Mux_v
    port map (
            O => \N__20300\,
            I => \N__20296\
        );

    \I__3463\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20293\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__20296\,
            I => \valueRegister_0_adj_1296\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__20293\,
            I => \valueRegister_0_adj_1296\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__3459\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20281\
        );

    \I__3458\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20278\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__20281\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__20278\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11\
        );

    \I__3455\ : InMux
    port map (
            O => \N__20273\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7924\
        );

    \I__3454\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20266\
        );

    \I__3453\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20263\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__20266\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__20263\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12\
        );

    \I__3450\ : InMux
    port map (
            O => \N__20258\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7925\
        );

    \I__3449\ : InMux
    port map (
            O => \N__20255\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7926\
        );

    \I__3448\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20248\
        );

    \I__3447\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20245\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__20248\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__20245\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14\
        );

    \I__3444\ : InMux
    port map (
            O => \N__20240\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7927\
        );

    \I__3443\ : InMux
    port map (
            O => \N__20237\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7928\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__20234\,
            I => \N__20230\
        );

    \I__3441\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20227\
        );

    \I__3440\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20224\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__20227\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__20224\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15\
        );

    \I__3437\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__3435\ : Span4Mux_v
    port map (
            O => \N__20213\,
            I => \N__20206\
        );

    \I__3434\ : InMux
    port map (
            O => \N__20212\,
            I => \N__20201\
        );

    \I__3433\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20201\
        );

    \I__3432\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20198\
        );

    \I__3431\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20195\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__20206\,
            I => \Inst_eia232.Inst_receiver.n7_adj_1264\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__20201\,
            I => \Inst_eia232.Inst_receiver.n7_adj_1264\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__20198\,
            I => \Inst_eia232.Inst_receiver.n7_adj_1264\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__20195\,
            I => \Inst_eia232.Inst_receiver.n7_adj_1264\
        );

    \I__3426\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20178\
        );

    \I__3425\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20165\
        );

    \I__3424\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20165\
        );

    \I__3423\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20165\
        );

    \I__3422\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20165\
        );

    \I__3421\ : InMux
    port map (
            O => \N__20181\,
            I => \N__20165\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20159\
        );

    \I__3419\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20154\
        );

    \I__3418\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20154\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__20165\,
            I => \N__20151\
        );

    \I__3416\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20144\
        );

    \I__3415\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20144\
        );

    \I__3414\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20144\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__20159\,
            I => \Inst_eia232.Inst_receiver.n957\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__20154\,
            I => \Inst_eia232.Inst_receiver.n957\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__20151\,
            I => \Inst_eia232.Inst_receiver.n957\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__20144\,
            I => \Inst_eia232.Inst_receiver.n957\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__20135\,
            I => \N__20130\
        );

    \I__3408\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20123\
        );

    \I__3407\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20123\
        );

    \I__3406\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20116\
        );

    \I__3405\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20116\
        );

    \I__3404\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20116\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__20123\,
            I => \N__20110\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__20116\,
            I => \N__20110\
        );

    \I__3401\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20107\
        );

    \I__3400\ : Span4Mux_h
    port map (
            O => \N__20110\,
            I => \N__20104\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__20107\,
            I => \Inst_eia232.Inst_receiver.bytecount_0\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__20104\,
            I => \Inst_eia232.Inst_receiver.bytecount_0\
        );

    \I__3397\ : CEMux
    port map (
            O => \N__20099\,
            I => \N__20095\
        );

    \I__3396\ : CEMux
    port map (
            O => \N__20098\,
            I => \N__20092\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__20095\,
            I => \N__20088\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__20092\,
            I => \N__20085\
        );

    \I__3393\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20082\
        );

    \I__3392\ : Span4Mux_h
    port map (
            O => \N__20088\,
            I => \N__20079\
        );

    \I__3391\ : Span4Mux_s1_v
    port map (
            O => \N__20085\,
            I => \N__20076\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__20082\,
            I => \N__20073\
        );

    \I__3389\ : Span4Mux_v
    port map (
            O => \N__20079\,
            I => \N__20070\
        );

    \I__3388\ : Span4Mux_v
    port map (
            O => \N__20076\,
            I => \N__20065\
        );

    \I__3387\ : Span4Mux_h
    port map (
            O => \N__20073\,
            I => \N__20065\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__20070\,
            I => \Inst_eia232.Inst_receiver.n3557\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__20065\,
            I => \Inst_eia232.Inst_receiver.n3557\
        );

    \I__3384\ : SRMux
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__20057\,
            I => \Inst_eia232.Inst_receiver.n8376\
        );

    \I__3382\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20050\
        );

    \I__3381\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20047\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__20050\,
            I => \configRegister_3_adj_1397\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__20047\,
            I => \configRegister_3_adj_1397\
        );

    \I__3378\ : InMux
    port map (
            O => \N__20042\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7916\
        );

    \I__3377\ : InMux
    port map (
            O => \N__20039\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7917\
        );

    \I__3376\ : InMux
    port map (
            O => \N__20036\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7918\
        );

    \I__3375\ : InMux
    port map (
            O => \N__20033\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7919\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__20030\,
            I => \N__20026\
        );

    \I__3373\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20023\
        );

    \I__3372\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20020\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__20023\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__20020\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7\
        );

    \I__3369\ : InMux
    port map (
            O => \N__20015\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7920\
        );

    \I__3368\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20008\
        );

    \I__3367\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20005\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__20005\,
            I => \configRegister_8_adj_1392\
        );

    \I__3364\ : Odrv12
    port map (
            O => \N__20002\,
            I => \configRegister_8_adj_1392\
        );

    \I__3363\ : InMux
    port map (
            O => \N__19997\,
            I => \bfn_6_4_0_\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__3361\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19987\
        );

    \I__3360\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__19987\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__19984\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9\
        );

    \I__3357\ : InMux
    port map (
            O => \N__19979\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7922\
        );

    \I__3356\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19972\
        );

    \I__3355\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19969\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__19972\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__19969\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10\
        );

    \I__3352\ : InMux
    port map (
            O => \N__19964\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7923\
        );

    \I__3351\ : InMux
    port map (
            O => \N__19961\,
            I => \bfn_6_3_0_\
        );

    \I__3350\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19954\
        );

    \I__3349\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19951\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__19954\,
            I => \configRegister_1_adj_1399\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__19951\,
            I => \configRegister_1_adj_1399\
        );

    \I__3346\ : InMux
    port map (
            O => \N__19946\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7914\
        );

    \I__3345\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__19940\,
            I => \N__19936\
        );

    \I__3343\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19933\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__19936\,
            I => \configRegister_2_adj_1398\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__19933\,
            I => \configRegister_2_adj_1398\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__3339\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19921\
        );

    \I__3338\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19918\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__19921\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__19918\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2\
        );

    \I__3335\ : InMux
    port map (
            O => \N__19913\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7915\
        );

    \I__3334\ : IoInMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__3332\ : Span4Mux_s0_v
    port map (
            O => \N__19904\,
            I => \N__19900\
        );

    \I__3331\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19897\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__19900\,
            I => testcnt_c_1
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__19897\,
            I => testcnt_c_1
        );

    \I__3328\ : InMux
    port map (
            O => \N__19892\,
            I => n7862
        );

    \I__3327\ : IoInMux
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__3325\ : IoSpan4Mux
    port map (
            O => \N__19883\,
            I => \N__19879\
        );

    \I__3324\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19876\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__19879\,
            I => testcnt_c_2
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__19876\,
            I => testcnt_c_2
        );

    \I__3321\ : InMux
    port map (
            O => \N__19871\,
            I => n7863
        );

    \I__3320\ : IoInMux
    port map (
            O => \N__19868\,
            I => \N__19864\
        );

    \I__3319\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19861\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__19864\,
            I => testcnt_c_3
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__19861\,
            I => testcnt_c_3
        );

    \I__3316\ : InMux
    port map (
            O => \N__19856\,
            I => n7864
        );

    \I__3315\ : IoInMux
    port map (
            O => \N__19853\,
            I => \N__19849\
        );

    \I__3314\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19846\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__19849\,
            I => testcnt_c_4
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__19846\,
            I => testcnt_c_4
        );

    \I__3311\ : InMux
    port map (
            O => \N__19841\,
            I => n7865
        );

    \I__3310\ : IoInMux
    port map (
            O => \N__19838\,
            I => \N__19834\
        );

    \I__3309\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__19834\,
            I => testcnt_c_5
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__19831\,
            I => testcnt_c_5
        );

    \I__3306\ : InMux
    port map (
            O => \N__19826\,
            I => n7866
        );

    \I__3305\ : IoInMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__3303\ : Span4Mux_s0_v
    port map (
            O => \N__19817\,
            I => \N__19813\
        );

    \I__3302\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19810\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__19813\,
            I => testcnt_c_6
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__19810\,
            I => testcnt_c_6
        );

    \I__3299\ : InMux
    port map (
            O => \N__19805\,
            I => n7867
        );

    \I__3298\ : InMux
    port map (
            O => \N__19802\,
            I => n7868
        );

    \I__3297\ : IoInMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__3295\ : Span4Mux_s0_v
    port map (
            O => \N__19793\,
            I => \N__19789\
        );

    \I__3294\ : InMux
    port map (
            O => \N__19792\,
            I => \N__19786\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__19789\,
            I => testcnt_c_7
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__19786\,
            I => testcnt_c_7
        );

    \I__3291\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__3289\ : Span4Mux_s2_v
    port map (
            O => \N__19775\,
            I => \N__19771\
        );

    \I__3288\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19768\
        );

    \I__3287\ : Span4Mux_v
    port map (
            O => \N__19771\,
            I => \N__19763\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__19768\,
            I => \N__19763\
        );

    \I__3285\ : Span4Mux_h
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__19760\,
            I => \GENERIC_FIFO_1.n8819\
        );

    \I__3283\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19753\
        );

    \I__3282\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19749\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__19753\,
            I => \N__19746\
        );

    \I__3280\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19742\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__19749\,
            I => \N__19736\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__19746\,
            I => \N__19736\
        );

    \I__3277\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19733\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19730\
        );

    \I__3275\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19726\
        );

    \I__3274\ : Span4Mux_v
    port map (
            O => \N__19736\,
            I => \N__19721\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__19733\,
            I => \N__19721\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__19730\,
            I => \N__19718\
        );

    \I__3271\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19715\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__19726\,
            I => \GENERIC_FIFO_1.read_pointer_7\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__19721\,
            I => \GENERIC_FIFO_1.read_pointer_7\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__19718\,
            I => \GENERIC_FIFO_1.read_pointer_7\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__19715\,
            I => \GENERIC_FIFO_1.read_pointer_7\
        );

    \I__3266\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19701\
        );

    \I__3265\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19695\
        );

    \I__3264\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19695\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__19701\,
            I => \N__19692\
        );

    \I__3262\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19679\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__19695\,
            I => \N__19676\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__19692\,
            I => \N__19673\
        );

    \I__3259\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19668\
        );

    \I__3258\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19668\
        );

    \I__3257\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19649\
        );

    \I__3256\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19649\
        );

    \I__3255\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19649\
        );

    \I__3254\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19649\
        );

    \I__3253\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19649\
        );

    \I__3252\ : InMux
    port map (
            O => \N__19684\,
            I => \N__19649\
        );

    \I__3251\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19649\
        );

    \I__3250\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19646\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19641\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__19676\,
            I => \N__19641\
        );

    \I__3247\ : Span4Mux_v
    port map (
            O => \N__19673\,
            I => \N__19636\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__19668\,
            I => \N__19636\
        );

    \I__3245\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19627\
        );

    \I__3244\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19627\
        );

    \I__3243\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19627\
        );

    \I__3242\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19627\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__19649\,
            I => \N__19624\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19619\
        );

    \I__3239\ : IoSpan4Mux
    port map (
            O => \N__19641\,
            I => \N__19619\
        );

    \I__3238\ : Span4Mux_h
    port map (
            O => \N__19636\,
            I => \N__19616\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__19627\,
            I => \N__19613\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__19624\,
            I => \N__19605\
        );

    \I__3235\ : Span4Mux_s1_v
    port map (
            O => \N__19619\,
            I => \N__19605\
        );

    \I__3234\ : Span4Mux_v
    port map (
            O => \N__19616\,
            I => \N__19605\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__19613\,
            I => \N__19602\
        );

    \I__3232\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19599\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__19605\,
            I => \GENERIC_FIFO_1.n141\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__19602\,
            I => \GENERIC_FIFO_1.n141\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__19599\,
            I => \GENERIC_FIFO_1.n141\
        );

    \I__3228\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__19589\,
            I => \N__19585\
        );

    \I__3226\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19582\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__19585\,
            I => \N__19579\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__19582\,
            I => \N__19576\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__19579\,
            I => \N__19573\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__19576\,
            I => \N__19570\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__19573\,
            I => \GENERIC_FIFO_1.n8820\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__19570\,
            I => \GENERIC_FIFO_1.n8820\
        );

    \I__3219\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19560\
        );

    \I__3218\ : InMux
    port map (
            O => \N__19564\,
            I => \N__19557\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__19563\,
            I => \N__19554\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__19560\,
            I => \N__19550\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__19557\,
            I => \N__19547\
        );

    \I__3214\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19544\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__19553\,
            I => \N__19541\
        );

    \I__3212\ : Span12Mux_v
    port map (
            O => \N__19550\,
            I => \N__19536\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__19547\,
            I => \N__19531\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19531\
        );

    \I__3209\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19526\
        );

    \I__3208\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19526\
        );

    \I__3207\ : InMux
    port map (
            O => \N__19539\,
            I => \N__19523\
        );

    \I__3206\ : Odrv12
    port map (
            O => \N__19536\,
            I => \GENERIC_FIFO_1.read_pointer_8\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__19531\,
            I => \GENERIC_FIFO_1.read_pointer_8\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__19526\,
            I => \GENERIC_FIFO_1.read_pointer_8\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__19523\,
            I => \GENERIC_FIFO_1.read_pointer_8\
        );

    \I__3202\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__3200\ : Odrv12
    port map (
            O => \N__19508\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_0\
        );

    \I__3199\ : SRMux
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__3197\ : Span4Mux_h
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__19496\,
            I => \Inst_core.Inst_sync.Inst_filter.n4732\
        );

    \I__3195\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__19490\,
            I => \Inst_core.Inst_sync.Inst_filter.input180Delay_4\
        );

    \I__3193\ : IoInMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__3191\ : Span4Mux_s0_v
    port map (
            O => \N__19481\,
            I => \N__19477\
        );

    \I__3190\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__19477\,
            I => testcnt_c_0
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__19474\,
            I => testcnt_c_0
        );

    \I__3187\ : InMux
    port map (
            O => \N__19469\,
            I => \bfn_6_1_0_\
        );

    \I__3186\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__3184\ : Span4Mux_h
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__19457\,
            I => \GENERIC_FIFO_1.n1424\
        );

    \I__3182\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__3180\ : Span4Mux_h
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__19445\,
            I => \GENERIC_FIFO_1.n1419\
        );

    \I__3178\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__19439\,
            I => \N__19435\
        );

    \I__3176\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__3175\ : Span4Mux_v
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__3173\ : Span4Mux_v
    port map (
            O => \N__19429\,
            I => \N__19423\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__19423\,
            I => \GENERIC_FIFO_1.n8813\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__19420\,
            I => \GENERIC_FIFO_1.n8813\
        );

    \I__3169\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19410\
        );

    \I__3168\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19407\
        );

    \I__3167\ : InMux
    port map (
            O => \N__19413\,
            I => \N__19404\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__19410\,
            I => \N__19401\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19397\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19392\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__19401\,
            I => \N__19392\
        );

    \I__3162\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19387\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__19397\,
            I => \N__19384\
        );

    \I__3160\ : Span4Mux_v
    port map (
            O => \N__19392\,
            I => \N__19381\
        );

    \I__3159\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19378\
        );

    \I__3158\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19375\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__19387\,
            I => \GENERIC_FIFO_1.read_pointer_1\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__19384\,
            I => \GENERIC_FIFO_1.read_pointer_1\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__19381\,
            I => \GENERIC_FIFO_1.read_pointer_1\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__19378\,
            I => \GENERIC_FIFO_1.read_pointer_1\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__19375\,
            I => \GENERIC_FIFO_1.read_pointer_1\
        );

    \I__3152\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__19361\,
            I => \N__19357\
        );

    \I__3150\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__3149\ : Span4Mux_v
    port map (
            O => \N__19357\,
            I => \N__19349\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__19354\,
            I => \N__19349\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__19346\,
            I => \GENERIC_FIFO_1.n8814\
        );

    \I__3145\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19339\
        );

    \I__3144\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19336\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__19339\,
            I => \N__19333\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__19336\,
            I => \N__19325\
        );

    \I__3141\ : Span4Mux_h
    port map (
            O => \N__19333\,
            I => \N__19325\
        );

    \I__3140\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19320\
        );

    \I__3139\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19320\
        );

    \I__3138\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19316\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__19325\,
            I => \N__19313\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__19320\,
            I => \N__19310\
        );

    \I__3135\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19307\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__19316\,
            I => \GENERIC_FIFO_1.read_pointer_2\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__19313\,
            I => \GENERIC_FIFO_1.read_pointer_2\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__19310\,
            I => \GENERIC_FIFO_1.read_pointer_2\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__19307\,
            I => \GENERIC_FIFO_1.read_pointer_2\
        );

    \I__3130\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__3128\ : Span4Mux_h
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__19289\,
            I => \GENERIC_FIFO_1.n1417\
        );

    \I__3126\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__19283\,
            I => \N__19279\
        );

    \I__3124\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19276\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__19279\,
            I => \N__19273\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__19276\,
            I => \N__19270\
        );

    \I__3121\ : Span4Mux_v
    port map (
            O => \N__19273\,
            I => \N__19267\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__19270\,
            I => \N__19264\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__19267\,
            I => \GENERIC_FIFO_1.n8816\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__19264\,
            I => \GENERIC_FIFO_1.n8816\
        );

    \I__3117\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19255\
        );

    \I__3116\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19252\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__19255\,
            I => \N__19249\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__19252\,
            I => \N__19241\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__19249\,
            I => \N__19241\
        );

    \I__3112\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19236\
        );

    \I__3111\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19236\
        );

    \I__3110\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19232\
        );

    \I__3109\ : Span4Mux_v
    port map (
            O => \N__19241\,
            I => \N__19227\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19227\
        );

    \I__3107\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19224\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__19232\,
            I => \GENERIC_FIFO_1.read_pointer_4\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__19227\,
            I => \GENERIC_FIFO_1.read_pointer_4\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__19224\,
            I => \GENERIC_FIFO_1.read_pointer_4\
        );

    \I__3103\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__19214\,
            I => \N__19210\
        );

    \I__3101\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19207\
        );

    \I__3100\ : Span4Mux_v
    port map (
            O => \N__19210\,
            I => \N__19204\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19201\
        );

    \I__3098\ : Span4Mux_h
    port map (
            O => \N__19204\,
            I => \N__19196\
        );

    \I__3097\ : Span4Mux_h
    port map (
            O => \N__19201\,
            I => \N__19196\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__19193\,
            I => \GENERIC_FIFO_1.n8817\
        );

    \I__3094\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__19187\,
            I => \N__19183\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__19186\,
            I => \N__19179\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__19183\,
            I => \N__19173\
        );

    \I__3090\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19170\
        );

    \I__3089\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19165\
        );

    \I__3088\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19165\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__19177\,
            I => \N__19162\
        );

    \I__3086\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19159\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__19173\,
            I => \N__19156\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__19170\,
            I => \N__19151\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19165\,
            I => \N__19151\
        );

    \I__3082\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19148\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__19159\,
            I => \GENERIC_FIFO_1.read_pointer_5\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__19156\,
            I => \GENERIC_FIFO_1.read_pointer_5\
        );

    \I__3079\ : Odrv4
    port map (
            O => \N__19151\,
            I => \GENERIC_FIFO_1.read_pointer_5\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__19148\,
            I => \GENERIC_FIFO_1.read_pointer_5\
        );

    \I__3077\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19132\
        );

    \I__3075\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19129\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__19132\,
            I => \N__19124\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__19129\,
            I => \N__19124\
        );

    \I__3072\ : Span4Mux_v
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__19121\,
            I => \GENERIC_FIFO_1.n8818\
        );

    \I__3070\ : InMux
    port map (
            O => \N__19118\,
            I => \N__19114\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__19117\,
            I => \N__19111\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19106\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19103\
        );

    \I__3066\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19100\
        );

    \I__3065\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19095\
        );

    \I__3064\ : Span12Mux_s4_h
    port map (
            O => \N__19106\,
            I => \N__19092\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__19103\,
            I => \N__19087\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__19100\,
            I => \N__19087\
        );

    \I__3061\ : InMux
    port map (
            O => \N__19099\,
            I => \N__19084\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19081\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__19095\,
            I => \GENERIC_FIFO_1.read_pointer_6\
        );

    \I__3058\ : Odrv12
    port map (
            O => \N__19092\,
            I => \GENERIC_FIFO_1.read_pointer_6\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__19087\,
            I => \GENERIC_FIFO_1.read_pointer_6\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__19084\,
            I => \GENERIC_FIFO_1.read_pointer_6\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__19081\,
            I => \GENERIC_FIFO_1.read_pointer_6\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__3053\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__3051\ : Span12Mux_s4_h
    port map (
            O => \N__19061\,
            I => \N__19057\
        );

    \I__3050\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19054\
        );

    \I__3049\ : Odrv12
    port map (
            O => \N__19057\,
            I => \valueRegister_4\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__19054\,
            I => \valueRegister_4\
        );

    \I__3047\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__19043\,
            I => \GENERIC_FIFO_1.n1422\
        );

    \I__3044\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__19037\,
            I => \N__19033\
        );

    \I__3042\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__19033\,
            I => \valueRegister_7\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__19030\,
            I => \valueRegister_7\
        );

    \I__3039\ : SRMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__3036\ : Span4Mux_s1_v
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__19013\,
            I => \Inst_core.Inst_sync.Inst_filter.n4729\
        );

    \I__3034\ : InMux
    port map (
            O => \N__19010\,
            I => \N__19007\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__19007\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_4\
        );

    \I__3032\ : InMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__19001\,
            I => \N__18997\
        );

    \I__3030\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18994\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__18997\,
            I => \N__18989\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__18994\,
            I => \N__18989\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__18989\,
            I => \N__18986\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__18983\,
            I => \GENERIC_FIFO_1.n8815\
        );

    \I__3024\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18976\
        );

    \I__3023\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18973\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18970\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__18973\,
            I => \N__18964\
        );

    \I__3020\ : Span4Mux_h
    port map (
            O => \N__18970\,
            I => \N__18964\
        );

    \I__3019\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18958\
        );

    \I__3018\ : Span4Mux_v
    port map (
            O => \N__18964\,
            I => \N__18955\
        );

    \I__3017\ : InMux
    port map (
            O => \N__18963\,
            I => \N__18952\
        );

    \I__3016\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18949\
        );

    \I__3015\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18946\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__18958\,
            I => \GENERIC_FIFO_1.read_pointer_3\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__18955\,
            I => \GENERIC_FIFO_1.read_pointer_3\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__18952\,
            I => \GENERIC_FIFO_1.read_pointer_3\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__18949\,
            I => \GENERIC_FIFO_1.read_pointer_3\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__18946\,
            I => \GENERIC_FIFO_1.read_pointer_3\
        );

    \I__3009\ : SRMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__3007\ : Span12Mux_s6_v
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__3006\ : Odrv12
    port map (
            O => \N__18926\,
            I => \Inst_core.Inst_sync.Inst_filter.n4731\
        );

    \I__3005\ : InMux
    port map (
            O => \N__18923\,
            I => \N__18919\
        );

    \I__3004\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18916\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__18919\,
            I => \maskRegister_2\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__18916\,
            I => \maskRegister_2\
        );

    \I__3001\ : SRMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__18899\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4740\
        );

    \I__2996\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18892\
        );

    \I__2995\ : InMux
    port map (
            O => \N__18895\,
            I => \N__18889\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__18892\,
            I => \N__18886\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__18889\,
            I => \maskRegister_3\
        );

    \I__2992\ : Odrv12
    port map (
            O => \N__18886\,
            I => \maskRegister_3\
        );

    \I__2991\ : SRMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__2989\ : Odrv12
    port map (
            O => \N__18875\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4741\
        );

    \I__2988\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18868\
        );

    \I__2987\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18865\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__18868\,
            I => \maskRegister_4\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__18865\,
            I => \maskRegister_4\
        );

    \I__2984\ : SRMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__2982\ : Span4Mux_h
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__18851\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4742\
        );

    \I__2980\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18844\
        );

    \I__2979\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18841\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__18844\,
            I => \maskRegister_6\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__18841\,
            I => \maskRegister_6\
        );

    \I__2976\ : SRMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__2974\ : Span4Mux_v
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__18827\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4744\
        );

    \I__2972\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18820\
        );

    \I__2971\ : InMux
    port map (
            O => \N__18823\,
            I => \N__18817\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__18820\,
            I => \maskRegister_7\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__18817\,
            I => \maskRegister_7\
        );

    \I__2968\ : SRMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__2966\ : Span4Mux_h
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__18803\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4745\
        );

    \I__2964\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18794\
        );

    \I__2963\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18794\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__18794\,
            I => \maskRegister_0_adj_1288\
        );

    \I__2961\ : SRMux
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__2959\ : Span4Mux_v
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__2958\ : Span4Mux_s1_h
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__18776\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4642\
        );

    \I__2955\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__18770\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_1\
        );

    \I__2953\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__18761\,
            I => \Inst_core.Inst_sync.Inst_filter.input360_2\
        );

    \I__2950\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__2948\ : Span12Mux_s4_h
    port map (
            O => \N__18752\,
            I => \N__18748\
        );

    \I__2947\ : InMux
    port map (
            O => \N__18751\,
            I => \N__18745\
        );

    \I__2946\ : Odrv12
    port map (
            O => \N__18748\,
            I => \valueRegister_6\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__18745\,
            I => \valueRegister_6\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_cascade_\
        );

    \I__2943\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18730\
        );

    \I__2942\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18730\
        );

    \I__2941\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18727\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__18730\,
            I => \N__18724\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__18727\,
            I => \configRegister_23_adj_1339\
        );

    \I__2938\ : Odrv12
    port map (
            O => \N__18724\,
            I => \configRegister_23_adj_1339\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__18719\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9090_cascade_\
        );

    \I__2936\ : SRMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18710\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__18710\,
            I => \Inst_core.Inst_sync.Inst_filter.n4730\
        );

    \I__2933\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18703\
        );

    \I__2932\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__18703\,
            I => \valueRegister_2\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__18700\,
            I => \valueRegister_2\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__2928\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18688\
        );

    \I__2927\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18685\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__18688\,
            I => \N__18682\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__18685\,
            I => \valueRegister_5\
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__18682\,
            I => \valueRegister_5\
        );

    \I__2923\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18673\
        );

    \I__2922\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18670\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__18673\,
            I => \configRegister_24\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__18670\,
            I => \configRegister_24\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__18665\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9096_cascade_\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__18662\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_cascade_\
        );

    \I__2917\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18654\
        );

    \I__2916\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18649\
        );

    \I__2915\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18649\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__18654\,
            I => \configRegister_23_adj_1379\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__18649\,
            I => \configRegister_23_adj_1379\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__18644\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9102_cascade_\
        );

    \I__2911\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18637\
        );

    \I__2910\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18634\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__18637\,
            I => \valueRegister_3\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__18634\,
            I => \valueRegister_3\
        );

    \I__2907\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18624\
        );

    \I__2906\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18619\
        );

    \I__2905\ : InMux
    port map (
            O => \N__18627\,
            I => \N__18619\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__18624\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__18619\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__18614\,
            I => \N__18611\
        );

    \I__2901\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18608\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__18608\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_3\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__18605\,
            I => \N__18601\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__18604\,
            I => \N__18598\
        );

    \I__2897\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18594\
        );

    \I__2896\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18589\
        );

    \I__2895\ : InMux
    port map (
            O => \N__18597\,
            I => \N__18589\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__18594\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__18589\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2\
        );

    \I__2892\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__18581\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_2\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__18578\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_cascade_\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__18575\,
            I => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9084_cascade_\
        );

    \I__2888\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__18569\,
            I => \N__18565\
        );

    \I__2886\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18562\
        );

    \I__2885\ : Span4Mux_v
    port map (
            O => \N__18565\,
            I => \N__18557\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__18562\,
            I => \N__18557\
        );

    \I__2883\ : Span4Mux_h
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__18554\,
            I => \N__18550\
        );

    \I__2881\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18547\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__18550\,
            I => \N__18544\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__18547\,
            I => \Inst_eia232.Inst_prescaler.counter_1\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__18544\,
            I => \Inst_eia232.Inst_prescaler.counter_1\
        );

    \I__2877\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18532\
        );

    \I__2875\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18529\
        );

    \I__2874\ : Span4Mux_h
    port map (
            O => \N__18532\,
            I => \N__18524\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__18529\,
            I => \N__18521\
        );

    \I__2872\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18516\
        );

    \I__2871\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18516\
        );

    \I__2870\ : Sp12to4
    port map (
            O => \N__18524\,
            I => \N__18511\
        );

    \I__2869\ : Span12Mux_s10_h
    port map (
            O => \N__18521\,
            I => \N__18511\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__18516\,
            I => \Inst_eia232.Inst_prescaler.counter_0\
        );

    \I__2867\ : Odrv12
    port map (
            O => \N__18511\,
            I => \Inst_eia232.Inst_prescaler.counter_0\
        );

    \I__2866\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18502\
        );

    \I__2865\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18499\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__18502\,
            I => \N__18496\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__18499\,
            I => \N__18493\
        );

    \I__2862\ : Odrv12
    port map (
            O => \N__18496\,
            I => \trxClock\
        );

    \I__2861\ : Odrv12
    port map (
            O => \N__18493\,
            I => \trxClock\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__2859\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18481\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__18484\,
            I => \N__18478\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__18481\,
            I => \N__18475\
        );

    \I__2856\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18472\
        );

    \I__2855\ : Span4Mux_s2_v
    port map (
            O => \N__18475\,
            I => \N__18465\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__18472\,
            I => \N__18465\
        );

    \I__2853\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18462\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__18470\,
            I => \N__18459\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__18465\,
            I => \N__18454\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__18462\,
            I => \N__18454\
        );

    \I__2849\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18451\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__18454\,
            I => \N__18446\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__18451\,
            I => \N__18446\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__2845\ : Span4Mux_v
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__18440\,
            I => \nstate_2__N_139_c_1\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_cascade_\
        );

    \I__2842\ : SRMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__2840\ : Span4Mux_s3_v
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__2839\ : Span4Mux_v
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__2838\ : Span4Mux_v
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__18419\,
            I => \Inst_eia232.Inst_prescaler.counter_4__N_38\
        );

    \I__2836\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18409\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__18415\,
            I => \N__18405\
        );

    \I__2834\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18400\
        );

    \I__2833\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18400\
        );

    \I__2832\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18397\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__18409\,
            I => \N__18394\
        );

    \I__2830\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18389\
        );

    \I__2829\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18389\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__18400\,
            I => \Inst_eia232.Inst_receiver.cmd_4\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__18397\,
            I => \Inst_eia232.Inst_receiver.cmd_4\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__18394\,
            I => \Inst_eia232.Inst_receiver.cmd_4\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__18389\,
            I => \Inst_eia232.Inst_receiver.cmd_4\
        );

    \I__2824\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__18377\,
            I => \N__18371\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__18376\,
            I => \N__18368\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__18375\,
            I => \N__18365\
        );

    \I__2820\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18360\
        );

    \I__2819\ : Span4Mux_h
    port map (
            O => \N__18371\,
            I => \N__18357\
        );

    \I__2818\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18348\
        );

    \I__2817\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18348\
        );

    \I__2816\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18348\
        );

    \I__2815\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18348\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__18360\,
            I => \Inst_eia232.Inst_receiver.cmd_5\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__18357\,
            I => \Inst_eia232.Inst_receiver.cmd_5\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__18348\,
            I => \Inst_eia232.Inst_receiver.cmd_5\
        );

    \I__2811\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18333\
        );

    \I__2810\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18333\
        );

    \I__2809\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18328\
        );

    \I__2808\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18328\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__18333\,
            I => n12
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__18328\,
            I => n12
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__2804\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18311\
        );

    \I__2803\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18311\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__18318\,
            I => \N__18304\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__18317\,
            I => \N__18299\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__18316\,
            I => \N__18296\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__18311\,
            I => \N__18290\
        );

    \I__2798\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18282\
        );

    \I__2797\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18282\
        );

    \I__2796\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18282\
        );

    \I__2795\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18279\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18274\
        );

    \I__2793\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18274\
        );

    \I__2792\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18261\
        );

    \I__2791\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18261\
        );

    \I__2790\ : InMux
    port map (
            O => \N__18296\,
            I => \N__18261\
        );

    \I__2789\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18261\
        );

    \I__2788\ : InMux
    port map (
            O => \N__18294\,
            I => \N__18261\
        );

    \I__2787\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18261\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__18290\,
            I => \N__18258\
        );

    \I__2785\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18255\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__18282\,
            I => \N__18252\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__18279\,
            I => \Inst_eia232.Inst_receiver.cmd_1\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__18274\,
            I => \Inst_eia232.Inst_receiver.cmd_1\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__18261\,
            I => \Inst_eia232.Inst_receiver.cmd_1\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__18258\,
            I => \Inst_eia232.Inst_receiver.cmd_1\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__18255\,
            I => \Inst_eia232.Inst_receiver.cmd_1\
        );

    \I__2778\ : Odrv4
    port map (
            O => \N__18252\,
            I => \Inst_eia232.Inst_receiver.cmd_1\
        );

    \I__2777\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18230\
        );

    \I__2776\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18230\
        );

    \I__2775\ : InMux
    port map (
            O => \N__18237\,
            I => \N__18230\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__18230\,
            I => \N__18222\
        );

    \I__2773\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18211\
        );

    \I__2772\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18211\
        );

    \I__2771\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18211\
        );

    \I__2770\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18211\
        );

    \I__2769\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18211\
        );

    \I__2768\ : Span4Mux_v
    port map (
            O => \N__18222\,
            I => \N__18208\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__18211\,
            I => \Inst_eia232.Inst_receiver.n3718\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__18208\,
            I => \Inst_eia232.Inst_receiver.n3718\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__18203\,
            I => \N__18195\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__18202\,
            I => \N__18190\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__18201\,
            I => \N__18186\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__18200\,
            I => \N__18183\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__18199\,
            I => \N__18180\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__18198\,
            I => \N__18174\
        );

    \I__2759\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18166\
        );

    \I__2758\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18166\
        );

    \I__2757\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18166\
        );

    \I__2756\ : InMux
    port map (
            O => \N__18190\,
            I => \N__18163\
        );

    \I__2755\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18148\
        );

    \I__2754\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18148\
        );

    \I__2753\ : InMux
    port map (
            O => \N__18183\,
            I => \N__18148\
        );

    \I__2752\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18148\
        );

    \I__2751\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18148\
        );

    \I__2750\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18148\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18148\
        );

    \I__2748\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18143\
        );

    \I__2747\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18143\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__18166\,
            I => \N__18140\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18163\,
            I => \Inst_eia232.Inst_receiver.cmd_2\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__18148\,
            I => \Inst_eia232.Inst_receiver.cmd_2\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__18143\,
            I => \Inst_eia232.Inst_receiver.cmd_2\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__18140\,
            I => \Inst_eia232.Inst_receiver.cmd_2\
        );

    \I__2741\ : InMux
    port map (
            O => \N__18131\,
            I => \N__18115\
        );

    \I__2740\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18115\
        );

    \I__2739\ : InMux
    port map (
            O => \N__18129\,
            I => \N__18115\
        );

    \I__2738\ : InMux
    port map (
            O => \N__18128\,
            I => \N__18098\
        );

    \I__2737\ : InMux
    port map (
            O => \N__18127\,
            I => \N__18098\
        );

    \I__2736\ : InMux
    port map (
            O => \N__18126\,
            I => \N__18098\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18098\
        );

    \I__2734\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18098\
        );

    \I__2733\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18098\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18098\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__18115\,
            I => \N__18095\
        );

    \I__2730\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18090\
        );

    \I__2729\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18090\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__18098\,
            I => \Inst_eia232.Inst_receiver.cmd_0\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__18095\,
            I => \Inst_eia232.Inst_receiver.cmd_0\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18090\,
            I => \Inst_eia232.Inst_receiver.cmd_0\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__18083\,
            I => \N__18076\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__18082\,
            I => \N__18070\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__18081\,
            I => \N__18066\
        );

    \I__2722\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18061\
        );

    \I__2721\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18061\
        );

    \I__2720\ : InMux
    port map (
            O => \N__18076\,
            I => \N__18042\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18075\,
            I => \N__18042\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18042\
        );

    \I__2717\ : InMux
    port map (
            O => \N__18073\,
            I => \N__18042\
        );

    \I__2716\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18042\
        );

    \I__2715\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18042\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18042\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__18061\,
            I => \N__18039\
        );

    \I__2712\ : InMux
    port map (
            O => \N__18060\,
            I => \N__18036\
        );

    \I__2711\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18029\
        );

    \I__2710\ : InMux
    port map (
            O => \N__18058\,
            I => \N__18029\
        );

    \I__2709\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18029\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__18042\,
            I => \N__18024\
        );

    \I__2707\ : Span4Mux_h
    port map (
            O => \N__18039\,
            I => \N__18024\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__18036\,
            I => \Inst_eia232.Inst_receiver.cmd_3\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__18029\,
            I => \Inst_eia232.Inst_receiver.cmd_3\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__18024\,
            I => \Inst_eia232.Inst_receiver.cmd_3\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__18017\,
            I => \N__18013\
        );

    \I__2702\ : InMux
    port map (
            O => \N__18016\,
            I => \N__18010\
        );

    \I__2701\ : InMux
    port map (
            O => \N__18013\,
            I => \N__18003\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__18010\,
            I => \N__18000\
        );

    \I__2699\ : InMux
    port map (
            O => \N__18009\,
            I => \N__17991\
        );

    \I__2698\ : InMux
    port map (
            O => \N__18008\,
            I => \N__17991\
        );

    \I__2697\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17991\
        );

    \I__2696\ : InMux
    port map (
            O => \N__18006\,
            I => \N__17991\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__18003\,
            I => \Inst_eia232.Inst_receiver.n69\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__18000\,
            I => \Inst_eia232.Inst_receiver.n69\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__17991\,
            I => \Inst_eia232.Inst_receiver.n69\
        );

    \I__2692\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17977\
        );

    \I__2691\ : InMux
    port map (
            O => \N__17983\,
            I => \N__17977\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__17982\,
            I => \N__17972\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__17977\,
            I => \N__17968\
        );

    \I__2688\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17962\
        );

    \I__2687\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17959\
        );

    \I__2686\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17954\
        );

    \I__2685\ : InMux
    port map (
            O => \N__17971\,
            I => \N__17954\
        );

    \I__2684\ : Span4Mux_h
    port map (
            O => \N__17968\,
            I => \N__17951\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__17967\,
            I => \N__17947\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__17966\,
            I => \N__17943\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__17965\,
            I => \N__17939\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__17962\,
            I => \N__17932\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__17959\,
            I => \N__17925\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__17954\,
            I => \N__17925\
        );

    \I__2677\ : Span4Mux_v
    port map (
            O => \N__17951\,
            I => \N__17925\
        );

    \I__2676\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17922\
        );

    \I__2675\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17911\
        );

    \I__2674\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17911\
        );

    \I__2673\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17911\
        );

    \I__2672\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17911\
        );

    \I__2671\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17911\
        );

    \I__2670\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17904\
        );

    \I__2669\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17904\
        );

    \I__2668\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17904\
        );

    \I__2667\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17901\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__17932\,
            I => \N__17896\
        );

    \I__2665\ : Span4Mux_v
    port map (
            O => \N__17925\,
            I => \N__17896\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__17922\,
            I => \Inst_eia232.state_1\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__17911\,
            I => \Inst_eia232.state_1\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__17904\,
            I => \Inst_eia232.state_1\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__17901\,
            I => \Inst_eia232.state_1\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__17896\,
            I => \Inst_eia232.state_1\
        );

    \I__2659\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17876\
        );

    \I__2658\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17876\
        );

    \I__2657\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17873\
        );

    \I__2656\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17870\
        );

    \I__2655\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17867\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__17876\,
            I => \N__17864\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17847\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__17870\,
            I => \N__17847\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17847\
        );

    \I__2650\ : Span4Mux_v
    port map (
            O => \N__17864\,
            I => \N__17847\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__17863\,
            I => \N__17843\
        );

    \I__2648\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17838\
        );

    \I__2647\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17835\
        );

    \I__2646\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17824\
        );

    \I__2645\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17824\
        );

    \I__2644\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17824\
        );

    \I__2643\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17824\
        );

    \I__2642\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17824\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__17847\,
            I => \N__17821\
        );

    \I__2640\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17812\
        );

    \I__2639\ : InMux
    port map (
            O => \N__17843\,
            I => \N__17812\
        );

    \I__2638\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17812\
        );

    \I__2637\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17812\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__17838\,
            I => \Inst_eia232.state_2\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__17835\,
            I => \Inst_eia232.state_2\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__17824\,
            I => \Inst_eia232.state_2\
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__17821\,
            I => \Inst_eia232.state_2\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__17812\,
            I => \Inst_eia232.state_2\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__17801\,
            I => \Inst_eia232.Inst_receiver.n7_cascade_\
        );

    \I__2630\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17788\
        );

    \I__2629\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17788\
        );

    \I__2628\ : InMux
    port map (
            O => \N__17796\,
            I => \N__17779\
        );

    \I__2627\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17779\
        );

    \I__2626\ : InMux
    port map (
            O => \N__17794\,
            I => \N__17779\
        );

    \I__2625\ : InMux
    port map (
            O => \N__17793\,
            I => \N__17779\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__17788\,
            I => \Inst_eia232.Inst_receiver.counter_1\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__17779\,
            I => \Inst_eia232.Inst_receiver.counter_1\
        );

    \I__2622\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17763\
        );

    \I__2621\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17763\
        );

    \I__2620\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17752\
        );

    \I__2619\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17752\
        );

    \I__2618\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17752\
        );

    \I__2617\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17752\
        );

    \I__2616\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17752\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__17763\,
            I => \Inst_eia232.Inst_receiver.counter_0\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__17752\,
            I => \Inst_eia232.Inst_receiver.counter_0\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__17747\,
            I => \N__17741\
        );

    \I__2612\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17735\
        );

    \I__2611\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17735\
        );

    \I__2610\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17728\
        );

    \I__2609\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17728\
        );

    \I__2608\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17728\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__17735\,
            I => \Inst_eia232.Inst_receiver.counter_2\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__17728\,
            I => \Inst_eia232.Inst_receiver.counter_2\
        );

    \I__2605\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17720\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__17720\,
            I => \Inst_eia232.Inst_receiver.n7777\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__17714\,
            I => \N__17711\
        );

    \I__2601\ : Span4Mux_s0_v
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__17708\,
            I => \Inst_eia232.Inst_receiver.n3202\
        );

    \I__2599\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17702\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__2597\ : Odrv12
    port map (
            O => \N__17699\,
            I => \Inst_eia232.Inst_receiver.n1_adj_1266\
        );

    \I__2596\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17687\
        );

    \I__2595\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17687\
        );

    \I__2594\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17680\
        );

    \I__2593\ : InMux
    port map (
            O => \N__17693\,
            I => \N__17680\
        );

    \I__2592\ : InMux
    port map (
            O => \N__17692\,
            I => \N__17680\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17677\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__17680\,
            I => \N__17668\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__17677\,
            I => \N__17668\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__17676\,
            I => \N__17665\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__17675\,
            I => \N__17658\
        );

    \I__2586\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17650\
        );

    \I__2585\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17647\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__17668\,
            I => \N__17644\
        );

    \I__2583\ : InMux
    port map (
            O => \N__17665\,
            I => \N__17633\
        );

    \I__2582\ : InMux
    port map (
            O => \N__17664\,
            I => \N__17633\
        );

    \I__2581\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17633\
        );

    \I__2580\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17633\
        );

    \I__2579\ : InMux
    port map (
            O => \N__17661\,
            I => \N__17633\
        );

    \I__2578\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17630\
        );

    \I__2577\ : InMux
    port map (
            O => \N__17657\,
            I => \N__17619\
        );

    \I__2576\ : InMux
    port map (
            O => \N__17656\,
            I => \N__17619\
        );

    \I__2575\ : InMux
    port map (
            O => \N__17655\,
            I => \N__17619\
        );

    \I__2574\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17619\
        );

    \I__2573\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17619\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__17650\,
            I => \Inst_eia232.state_0\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__17647\,
            I => \Inst_eia232.state_0\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__17644\,
            I => \Inst_eia232.state_0\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__17633\,
            I => \Inst_eia232.state_0\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__17630\,
            I => \Inst_eia232.state_0\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__17619\,
            I => \Inst_eia232.state_0\
        );

    \I__2566\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17599\
        );

    \I__2565\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17592\
        );

    \I__2564\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17592\
        );

    \I__2563\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17592\
        );

    \I__2562\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17589\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__17599\,
            I => \N__17584\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__17592\,
            I => \N__17584\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__17589\,
            I => \Inst_eia232.Inst_receiver.nstate_2_N_133_1\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__17584\,
            I => \Inst_eia232.Inst_receiver.nstate_2_N_133_1\
        );

    \I__2557\ : InMux
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__2555\ : Odrv12
    port map (
            O => \N__17573\,
            I => \Inst_eia232.Inst_receiver.n8826\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__17570\,
            I => \Inst_eia232.Inst_receiver.n3504_cascade_\
        );

    \I__2553\ : CEMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__17561\,
            I => \N__17558\
        );

    \I__2550\ : Span4Mux_s0_v
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__17555\,
            I => \Inst_eia232.Inst_receiver.n3676\
        );

    \I__2548\ : SRMux
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__17543\,
            I => \Inst_eia232.Inst_receiver.n4767\
        );

    \I__2544\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__17537\,
            I => \Inst_eia232.Inst_receiver.n3504\
        );

    \I__2542\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17528\
        );

    \I__2541\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17528\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__17525\,
            I => \Inst_eia232.Inst_receiver.n5\
        );

    \I__2538\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17515\
        );

    \I__2537\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17515\
        );

    \I__2536\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17512\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__17515\,
            I => \Inst_eia232.Inst_receiver.n75\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__17512\,
            I => \Inst_eia232.Inst_receiver.n75\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__17507\,
            I => \N__17504\
        );

    \I__2532\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17498\
        );

    \I__2531\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17498\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__17498\,
            I => \Inst_eia232.Inst_receiver.n14\
        );

    \I__2529\ : SRMux
    port map (
            O => \N__17495\,
            I => \N__17491\
        );

    \I__2528\ : SRMux
    port map (
            O => \N__17494\,
            I => \N__17488\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__17491\,
            I => \N__17483\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__17488\,
            I => \N__17480\
        );

    \I__2525\ : SRMux
    port map (
            O => \N__17487\,
            I => \N__17477\
        );

    \I__2524\ : SRMux
    port map (
            O => \N__17486\,
            I => \N__17474\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__17483\,
            I => \N__17471\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__17480\,
            I => \N__17464\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__17477\,
            I => \N__17464\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__17474\,
            I => \N__17464\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__17471\,
            I => n1917
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__17464\,
            I => n1917
        );

    \I__2517\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17449\
        );

    \I__2516\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17449\
        );

    \I__2515\ : InMux
    port map (
            O => \N__17457\,
            I => \N__17449\
        );

    \I__2514\ : InMux
    port map (
            O => \N__17456\,
            I => \N__17446\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__17449\,
            I => \Inst_eia232.Inst_receiver.counter_4\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__17446\,
            I => \Inst_eia232.Inst_receiver.counter_4\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__17441\,
            I => \N__17436\
        );

    \I__2510\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17431\
        );

    \I__2509\ : InMux
    port map (
            O => \N__17439\,
            I => \N__17428\
        );

    \I__2508\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17421\
        );

    \I__2507\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17421\
        );

    \I__2506\ : InMux
    port map (
            O => \N__17434\,
            I => \N__17421\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__17431\,
            I => \Inst_eia232.Inst_receiver.counter_3\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__17428\,
            I => \Inst_eia232.Inst_receiver.counter_3\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__17421\,
            I => \Inst_eia232.Inst_receiver.counter_3\
        );

    \I__2502\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17409\
        );

    \I__2501\ : InMux
    port map (
            O => \N__17413\,
            I => \N__17404\
        );

    \I__2500\ : InMux
    port map (
            O => \N__17412\,
            I => \N__17404\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__17409\,
            I => \Inst_eia232.Inst_receiver.n5504\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__17404\,
            I => \Inst_eia232.Inst_receiver.n5504\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__17399\,
            I => \Inst_eia232.Inst_receiver.n8782_cascade_\
        );

    \I__2496\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17390\
        );

    \I__2495\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17390\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__17390\,
            I => \Inst_eia232.Inst_receiver.n6_adj_1267\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__17387\,
            I => \Inst_eia232.Inst_receiver.n3_cascade_\
        );

    \I__2492\ : InMux
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__17381\,
            I => \Inst_eia232.Inst_receiver.n5505\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__17378\,
            I => \Inst_eia232.Inst_receiver.n8755_cascade_\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__17375\,
            I => \Inst_eia232.Inst_receiver.n9123_cascade_\
        );

    \I__2488\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__17369\,
            I => \executePrev\
        );

    \I__2486\ : InMux
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__17363\,
            I => \Inst_eia232.Inst_receiver.n8784\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__17360\,
            I => \Inst_eia232.Inst_receiver.n6_cascade_\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__17357\,
            I => \Inst_eia232.Inst_receiver.n8_cascade_\
        );

    \I__2482\ : SRMux
    port map (
            O => \N__17354\,
            I => \N__17351\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__17351\,
            I => \N__17346\
        );

    \I__2480\ : SRMux
    port map (
            O => \N__17350\,
            I => \N__17343\
        );

    \I__2479\ : InMux
    port map (
            O => \N__17349\,
            I => \N__17340\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__17346\,
            I => \N__17335\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__17343\,
            I => \N__17335\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17332\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__17335\,
            I => \N__17329\
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__17332\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__17329\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2472\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__17321\,
            I => \GENERIC_FIFO_1.n1388\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__17318\,
            I => \N__17315\
        );

    \I__2469\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17312\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__17312\,
            I => \N__17309\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__17309\,
            I => \GENERIC_FIFO_1.n1373\
        );

    \I__2466\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17303\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__2464\ : Span4Mux_s3_h
    port map (
            O => \N__17300\,
            I => \N__17297\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__17297\,
            I => \N__17294\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__17294\,
            I => \GENERIC_FIFO_1.n8630\
        );

    \I__2461\ : InMux
    port map (
            O => \N__17291\,
            I => \bfn_4_16_0_\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__17288\,
            I => \N__17285\
        );

    \I__2459\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17282\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__17279\,
            I => \GENERIC_FIFO_1.n1372\
        );

    \I__2456\ : InMux
    port map (
            O => \N__17276\,
            I => \GENERIC_FIFO_1.n7945\
        );

    \I__2455\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17270\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__17270\,
            I => \GENERIC_FIFO_1.n1383\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2452\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__17261\,
            I => \N__17258\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__17258\,
            I => \GENERIC_FIFO_1.n1371\
        );

    \I__2449\ : InMux
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__17252\,
            I => \N__17249\
        );

    \I__2447\ : Span4Mux_v
    port map (
            O => \N__17249\,
            I => \N__17246\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__17246\,
            I => \N__17243\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__17243\,
            I => \GENERIC_FIFO_1.n8638\
        );

    \I__2444\ : InMux
    port map (
            O => \N__17240\,
            I => \GENERIC_FIFO_1.n7946\
        );

    \I__2443\ : InMux
    port map (
            O => \N__17237\,
            I => \GENERIC_FIFO_1.n1392\
        );

    \I__2442\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17230\
        );

    \I__2441\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17226\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__17230\,
            I => \N__17223\
        );

    \I__2439\ : InMux
    port map (
            O => \N__17229\,
            I => \N__17220\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__17226\,
            I => \N__17217\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__17223\,
            I => \N__17212\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__17220\,
            I => \N__17212\
        );

    \I__2435\ : Span4Mux_s3_h
    port map (
            O => \N__17217\,
            I => \N__17209\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__17212\,
            I => \N__17206\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__17209\,
            I => \GENERIC_FIFO_1.n1392_THRU_CO\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__17206\,
            I => \GENERIC_FIFO_1.n1392_THRU_CO\
        );

    \I__2431\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__2429\ : Span4Mux_s3_v
    port map (
            O => \N__17195\,
            I => \N__17191\
        );

    \I__2428\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17188\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__17191\,
            I => \N__17185\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__17188\,
            I => \N__17182\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__17185\,
            I => \GENERIC_FIFO_1.n8821\
        );

    \I__2424\ : Odrv12
    port map (
            O => \N__17182\,
            I => \GENERIC_FIFO_1.n8821\
        );

    \I__2423\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17173\
        );

    \I__2422\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17169\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__17173\,
            I => \N__17166\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__17172\,
            I => \N__17163\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__17169\,
            I => \N__17158\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__17166\,
            I => \N__17158\
        );

    \I__2417\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17155\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__17158\,
            I => \N__17149\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__17155\,
            I => \N__17146\
        );

    \I__2414\ : InMux
    port map (
            O => \N__17154\,
            I => \N__17139\
        );

    \I__2413\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17139\
        );

    \I__2412\ : InMux
    port map (
            O => \N__17152\,
            I => \N__17139\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__17149\,
            I => \GENERIC_FIFO_1.read_pointer_9\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__17146\,
            I => \GENERIC_FIFO_1.read_pointer_9\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__17139\,
            I => \GENERIC_FIFO_1.read_pointer_9\
        );

    \I__2408\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__17129\,
            I => \N__17126\
        );

    \I__2406\ : Span4Mux_s3_h
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__17123\,
            I => \GENERIC_FIFO_1.n1416\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__2403\ : CascadeBuf
    port map (
            O => \N__17117\,
            I => \N__17112\
        );

    \I__2402\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17109\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17106\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__17112\,
            I => \N__17103\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17109\,
            I => \N__17098\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__17106\,
            I => \N__17095\
        );

    \I__2397\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17092\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17089\
        );

    \I__2395\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17086\
        );

    \I__2394\ : Span4Mux_s2_v
    port map (
            O => \N__17098\,
            I => \N__17081\
        );

    \I__2393\ : Span4Mux_h
    port map (
            O => \N__17095\,
            I => \N__17081\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__17092\,
            I => \N__17078\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__17089\,
            I => \GENERIC_FIFO_1.write_pointer_6\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__17086\,
            I => \GENERIC_FIFO_1.write_pointer_6\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__17081\,
            I => \GENERIC_FIFO_1.write_pointer_6\
        );

    \I__2388\ : Odrv12
    port map (
            O => \N__17078\,
            I => \GENERIC_FIFO_1.write_pointer_6\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17066\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__17066\,
            I => \N__17061\
        );

    \I__2385\ : InMux
    port map (
            O => \N__17065\,
            I => \N__17058\
        );

    \I__2384\ : InMux
    port map (
            O => \N__17064\,
            I => \N__17053\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__17061\,
            I => \N__17047\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__17058\,
            I => \N__17047\
        );

    \I__2381\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17044\
        );

    \I__2380\ : InMux
    port map (
            O => \N__17056\,
            I => \N__17041\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__17038\
        );

    \I__2378\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17035\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__17047\,
            I => \N__17030\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__17044\,
            I => \N__17030\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__17041\,
            I => \N__17025\
        );

    \I__2374\ : Span12Mux_s2_v
    port map (
            O => \N__17038\,
            I => \N__17025\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__17035\,
            I => \GENERIC_FIFO_1.read_pointer_0\
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__17030\,
            I => \GENERIC_FIFO_1.read_pointer_0\
        );

    \I__2371\ : Odrv12
    port map (
            O => \N__17025\,
            I => \GENERIC_FIFO_1.read_pointer_0\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__2369\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__17012\,
            I => \GENERIC_FIFO_1.n2\
        );

    \I__2367\ : InMux
    port map (
            O => \N__17009\,
            I => \bfn_4_15_0_\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__2365\ : InMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__17000\,
            I => \GENERIC_FIFO_1.n1379\
        );

    \I__2363\ : InMux
    port map (
            O => \N__16997\,
            I => \GENERIC_FIFO_1.n7938\
        );

    \I__2362\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__16991\,
            I => \GENERIC_FIFO_1.n1391\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__2359\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__2357\ : Odrv12
    port map (
            O => \N__16979\,
            I => \GENERIC_FIFO_1.n1378\
        );

    \I__2356\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__16973\,
            I => \N__16970\
        );

    \I__2354\ : Span4Mux_s3_h
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__16967\,
            I => \N__16964\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__16964\,
            I => \GENERIC_FIFO_1.n8634\
        );

    \I__2351\ : InMux
    port map (
            O => \N__16961\,
            I => \GENERIC_FIFO_1.n7939\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__2349\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__16952\,
            I => \GENERIC_FIFO_1.n1377\
        );

    \I__2347\ : InMux
    port map (
            O => \N__16949\,
            I => \GENERIC_FIFO_1.n7940\
        );

    \I__2346\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__16943\,
            I => \GENERIC_FIFO_1.n1390\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__16940\,
            I => \N__16937\
        );

    \I__2343\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__16928\,
            I => \GENERIC_FIFO_1.n1376\
        );

    \I__2339\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__16922\,
            I => \N__16919\
        );

    \I__2337\ : Span4Mux_s3_h
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__2336\ : Span4Mux_v
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__16913\,
            I => \GENERIC_FIFO_1.n8628\
        );

    \I__2334\ : InMux
    port map (
            O => \N__16910\,
            I => \GENERIC_FIFO_1.n7941\
        );

    \I__2333\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16904\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__2331\ : Span4Mux_s2_v
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__16898\,
            I => \GENERIC_FIFO_1.n1375\
        );

    \I__2329\ : InMux
    port map (
            O => \N__16895\,
            I => \GENERIC_FIFO_1.n7942\
        );

    \I__2328\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__16889\,
            I => \GENERIC_FIFO_1.n1386\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__2325\ : InMux
    port map (
            O => \N__16883\,
            I => \N__16880\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__16880\,
            I => \GENERIC_FIFO_1.n1374\
        );

    \I__2323\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16874\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__16874\,
            I => \N__16871\
        );

    \I__2321\ : Span12Mux_v
    port map (
            O => \N__16871\,
            I => \N__16868\
        );

    \I__2320\ : Odrv12
    port map (
            O => \N__16868\,
            I => \GENERIC_FIFO_1.n8632\
        );

    \I__2319\ : InMux
    port map (
            O => \N__16865\,
            I => \GENERIC_FIFO_1.n7943\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__16862\,
            I => \N__16859\
        );

    \I__2317\ : InMux
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__16856\,
            I => \N__16853\
        );

    \I__2315\ : Span4Mux_s3_h
    port map (
            O => \N__16853\,
            I => \N__16850\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__16850\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_7\
        );

    \I__2313\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__16844\,
            I => \GENERIC_FIFO_1.n17_adj_1280\
        );

    \I__2311\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__16835\,
            I => \GENERIC_FIFO_1.n1421\
        );

    \I__2308\ : InMux
    port map (
            O => \N__16832\,
            I => \N__16829\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__16829\,
            I => \N__16826\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__16826\,
            I => \GENERIC_FIFO_1.n1423\
        );

    \I__2305\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16819\
        );

    \I__2304\ : SRMux
    port map (
            O => \N__16822\,
            I => \N__16816\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__16819\,
            I => \N__16808\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__16816\,
            I => \N__16808\
        );

    \I__2301\ : SRMux
    port map (
            O => \N__16815\,
            I => \N__16805\
        );

    \I__2300\ : SRMux
    port map (
            O => \N__16814\,
            I => \N__16799\
        );

    \I__2299\ : InMux
    port map (
            O => \N__16813\,
            I => \N__16796\
        );

    \I__2298\ : Span4Mux_s3_v
    port map (
            O => \N__16808\,
            I => \N__16784\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__16805\,
            I => \N__16784\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__16804\,
            I => \N__16780\
        );

    \I__2295\ : InMux
    port map (
            O => \N__16803\,
            I => \N__16773\
        );

    \I__2294\ : InMux
    port map (
            O => \N__16802\,
            I => \N__16773\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__16799\,
            I => \N__16770\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__16796\,
            I => \N__16767\
        );

    \I__2291\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16752\
        );

    \I__2290\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16752\
        );

    \I__2289\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16752\
        );

    \I__2288\ : InMux
    port map (
            O => \N__16792\,
            I => \N__16752\
        );

    \I__2287\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16752\
        );

    \I__2286\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16752\
        );

    \I__2285\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16752\
        );

    \I__2284\ : Span4Mux_v
    port map (
            O => \N__16784\,
            I => \N__16749\
        );

    \I__2283\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16740\
        );

    \I__2282\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16740\
        );

    \I__2281\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16740\
        );

    \I__2280\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16740\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__16773\,
            I => \N__16737\
        );

    \I__2278\ : Sp12to4
    port map (
            O => \N__16770\,
            I => \N__16732\
        );

    \I__2277\ : Span12Mux_s11_h
    port map (
            O => \N__16767\,
            I => \N__16732\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__16752\,
            I => \writeByte\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__16749\,
            I => \writeByte\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__16740\,
            I => \writeByte\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__16737\,
            I => \writeByte\
        );

    \I__2272\ : Odrv12
    port map (
            O => \N__16732\,
            I => \writeByte\
        );

    \I__2271\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__16718\,
            I => \N__16714\
        );

    \I__2269\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16711\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__16714\,
            I => \N__16708\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__16711\,
            I => \N__16703\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__16708\,
            I => \N__16700\
        );

    \I__2265\ : InMux
    port map (
            O => \N__16707\,
            I => \N__16695\
        );

    \I__2264\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16695\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__16703\,
            I => n9
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__16700\,
            I => n9
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__16695\,
            I => n9
        );

    \I__2260\ : SRMux
    port map (
            O => \N__16688\,
            I => \N__16682\
        );

    \I__2259\ : SRMux
    port map (
            O => \N__16687\,
            I => \N__16679\
        );

    \I__2258\ : CEMux
    port map (
            O => \N__16686\,
            I => \N__16676\
        );

    \I__2257\ : CEMux
    port map (
            O => \N__16685\,
            I => \N__16673\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__16682\,
            I => \N__16670\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__16679\,
            I => \N__16667\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__16676\,
            I => \N__16664\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__16673\,
            I => \N__16661\
        );

    \I__2252\ : Span4Mux_s3_h
    port map (
            O => \N__16670\,
            I => \N__16658\
        );

    \I__2251\ : Span4Mux_s3_h
    port map (
            O => \N__16667\,
            I => \N__16655\
        );

    \I__2250\ : Span12Mux_s3_h
    port map (
            O => \N__16664\,
            I => \N__16652\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__16661\,
            I => \N__16649\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__16658\,
            I => \N__16646\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__16655\,
            I => \N__16643\
        );

    \I__2246\ : Odrv12
    port map (
            O => \N__16652\,
            I => \Inst_eia232.Inst_transmitter.n3608\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__16649\,
            I => \Inst_eia232.Inst_transmitter.n3608\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__16646\,
            I => \Inst_eia232.Inst_transmitter.n3608\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__16643\,
            I => \Inst_eia232.Inst_transmitter.n3608\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__16634\,
            I => \N__16631\
        );

    \I__2241\ : CascadeBuf
    port map (
            O => \N__16631\,
            I => \N__16626\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__16630\,
            I => \N__16623\
        );

    \I__2239\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16620\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__16626\,
            I => \N__16617\
        );

    \I__2237\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16612\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__16620\,
            I => \N__16609\
        );

    \I__2235\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16606\
        );

    \I__2234\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16603\
        );

    \I__2233\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16600\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__16612\,
            I => \N__16597\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__16609\,
            I => \N__16592\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__16606\,
            I => \N__16592\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__16603\,
            I => \GENERIC_FIFO_1.write_pointer_0\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__16600\,
            I => \GENERIC_FIFO_1.write_pointer_0\
        );

    \I__2227\ : Odrv12
    port map (
            O => \N__16597\,
            I => \GENERIC_FIFO_1.write_pointer_0\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__16592\,
            I => \GENERIC_FIFO_1.write_pointer_0\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__2224\ : CascadeBuf
    port map (
            O => \N__16580\,
            I => \N__16576\
        );

    \I__2223\ : InMux
    port map (
            O => \N__16579\,
            I => \N__16572\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__16576\,
            I => \N__16569\
        );

    \I__2221\ : InMux
    port map (
            O => \N__16575\,
            I => \N__16564\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__16572\,
            I => \N__16561\
        );

    \I__2219\ : InMux
    port map (
            O => \N__16569\,
            I => \N__16558\
        );

    \I__2218\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16555\
        );

    \I__2217\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16552\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__16564\,
            I => \N__16549\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__16561\,
            I => \N__16544\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__16558\,
            I => \N__16544\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__16555\,
            I => \GENERIC_FIFO_1.write_pointer_1\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__16552\,
            I => \GENERIC_FIFO_1.write_pointer_1\
        );

    \I__2211\ : Odrv12
    port map (
            O => \N__16549\,
            I => \GENERIC_FIFO_1.write_pointer_1\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__16544\,
            I => \GENERIC_FIFO_1.write_pointer_1\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__2208\ : CascadeBuf
    port map (
            O => \N__16532\,
            I => \N__16527\
        );

    \I__2207\ : InMux
    port map (
            O => \N__16531\,
            I => \N__16524\
        );

    \I__2206\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16521\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__16527\,
            I => \N__16518\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__16524\,
            I => \N__16513\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__16521\,
            I => \N__16510\
        );

    \I__2202\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16507\
        );

    \I__2201\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16504\
        );

    \I__2200\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16501\
        );

    \I__2199\ : Span4Mux_v
    port map (
            O => \N__16513\,
            I => \N__16494\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__16510\,
            I => \N__16494\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__16507\,
            I => \N__16494\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__16504\,
            I => \GENERIC_FIFO_1.write_pointer_2\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__16501\,
            I => \GENERIC_FIFO_1.write_pointer_2\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__16494\,
            I => \GENERIC_FIFO_1.write_pointer_2\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__2192\ : CascadeBuf
    port map (
            O => \N__16484\,
            I => \N__16479\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16483\,
            I => \N__16476\
        );

    \I__2190\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16473\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__16479\,
            I => \N__16470\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__16476\,
            I => \N__16465\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__16473\,
            I => \N__16462\
        );

    \I__2186\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16459\
        );

    \I__2185\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16456\
        );

    \I__2184\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16453\
        );

    \I__2183\ : Span4Mux_v
    port map (
            O => \N__16465\,
            I => \N__16446\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__16462\,
            I => \N__16446\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__16459\,
            I => \N__16446\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__16456\,
            I => \GENERIC_FIFO_1.write_pointer_3\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__16453\,
            I => \GENERIC_FIFO_1.write_pointer_3\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__16446\,
            I => \GENERIC_FIFO_1.write_pointer_3\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__2176\ : CascadeBuf
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16427\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__16427\,
            I => \GENERIC_FIFO_1.n76\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__16424\,
            I => \N__16421\
        );

    \I__2171\ : CascadeBuf
    port map (
            O => \N__16421\,
            I => \N__16418\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__16418\,
            I => \N__16415\
        );

    \I__2169\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__16412\,
            I => \GENERIC_FIFO_1.n75\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__2166\ : CascadeBuf
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__16403\,
            I => \N__16400\
        );

    \I__2164\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__16397\,
            I => \GENERIC_FIFO_1.n74\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__16394\,
            I => \N__16391\
        );

    \I__2161\ : CascadeBuf
    port map (
            O => \N__16391\,
            I => \N__16388\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__2159\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__16382\,
            I => \GENERIC_FIFO_1.n73\
        );

    \I__2157\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16376\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__16376\,
            I => \N__16373\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__16370\,
            I => \GENERIC_FIFO_1.n1420\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__16367\,
            I => \N__16364\
        );

    \I__2152\ : CascadeBuf
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__2150\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16355\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__16355\,
            I => \GENERIC_FIFO_1.n72\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__16352\,
            I => \GENERIC_FIFO_1.n16_adj_1279_cascade_\
        );

    \I__2147\ : InMux
    port map (
            O => \N__16349\,
            I => \N__16331\
        );

    \I__2146\ : InMux
    port map (
            O => \N__16348\,
            I => \N__16331\
        );

    \I__2145\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16331\
        );

    \I__2144\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16331\
        );

    \I__2143\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16328\
        );

    \I__2142\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16325\
        );

    \I__2141\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16316\
        );

    \I__2140\ : InMux
    port map (
            O => \N__16342\,
            I => \N__16316\
        );

    \I__2139\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16316\
        );

    \I__2138\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16316\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__16331\,
            I => \N__16313\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__16328\,
            I => \N__16308\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__16325\,
            I => \N__16308\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__16316\,
            I => \N__16305\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__16313\,
            I => \N__16302\
        );

    \I__2132\ : Span4Mux_s2_h
    port map (
            O => \N__16308\,
            I => \N__16297\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__16305\,
            I => \N__16297\
        );

    \I__2130\ : Span4Mux_v
    port map (
            O => \N__16302\,
            I => \N__16292\
        );

    \I__2129\ : Span4Mux_v
    port map (
            O => \N__16297\,
            I => \N__16292\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__16292\,
            I => \GENERIC_FIFO_1.n142\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__16289\,
            I => \N__16286\
        );

    \I__2126\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16283\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__16283\,
            I => \N__16280\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__16280\,
            I => \N__16277\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__16277\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_7\
        );

    \I__2122\ : SRMux
    port map (
            O => \N__16274\,
            I => \N__16271\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__16271\,
            I => \N__16268\
        );

    \I__2120\ : Span4Mux_s2_v
    port map (
            O => \N__16268\,
            I => \N__16265\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__16265\,
            I => \N__16262\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__16262\,
            I => \Inst_eia232.Inst_receiver.n4628\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16256\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__16256\,
            I => \N__16253\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__16253\,
            I => \N__16250\
        );

    \I__2114\ : Span4Mux_h
    port map (
            O => \N__16250\,
            I => \N__16246\
        );

    \I__2113\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16243\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__16246\,
            I => \N__16238\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__16243\,
            I => \N__16238\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__16238\,
            I => \N__16235\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__16235\,
            I => \Inst_eia232.Inst_transmitter.paused\
        );

    \I__2108\ : SRMux
    port map (
            O => \N__16232\,
            I => \N__16229\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__16229\,
            I => \N__16225\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__16228\,
            I => \N__16222\
        );

    \I__2105\ : Span4Mux_s2_h
    port map (
            O => \N__16225\,
            I => \N__16217\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__16222\,
            I => \N__16217\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__16217\,
            I => \N__16214\
        );

    \I__2102\ : Span4Mux_v
    port map (
            O => \N__16214\,
            I => \N__16211\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__16211\,
            I => \Inst_eia232.Inst_transmitter.n4634\
        );

    \I__2100\ : SRMux
    port map (
            O => \N__16208\,
            I => \N__16199\
        );

    \I__2099\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16199\
        );

    \I__2098\ : InMux
    port map (
            O => \N__16206\,
            I => \N__16199\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__16199\,
            I => \N__16193\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__16198\,
            I => \N__16188\
        );

    \I__2095\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16182\
        );

    \I__2094\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16182\
        );

    \I__2093\ : Span4Mux_h
    port map (
            O => \N__16193\,
            I => \N__16179\
        );

    \I__2092\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16174\
        );

    \I__2091\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16170\
        );

    \I__2090\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16165\
        );

    \I__2089\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16165\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__16182\,
            I => \N__16160\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__16179\,
            I => \N__16160\
        );

    \I__2086\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16155\
        );

    \I__2085\ : InMux
    port map (
            O => \N__16177\,
            I => \N__16155\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__16174\,
            I => \N__16152\
        );

    \I__2083\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16149\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__16170\,
            I => state_0
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__16165\,
            I => state_0
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__16160\,
            I => state_0
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__16155\,
            I => state_0
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__16152\,
            I => state_0
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__16149\,
            I => state_0
        );

    \I__2076\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16133\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__16133\,
            I => \N__16125\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__16132\,
            I => \N__16122\
        );

    \I__2073\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16112\
        );

    \I__2072\ : InMux
    port map (
            O => \N__16130\,
            I => \N__16112\
        );

    \I__2071\ : InMux
    port map (
            O => \N__16129\,
            I => \N__16112\
        );

    \I__2070\ : InMux
    port map (
            O => \N__16128\,
            I => \N__16112\
        );

    \I__2069\ : Span4Mux_h
    port map (
            O => \N__16125\,
            I => \N__16109\
        );

    \I__2068\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16104\
        );

    \I__2067\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16104\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__16112\,
            I => \N__16101\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__16109\,
            I => \N__16098\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__16104\,
            I => \Inst_eia232.Inst_transmitter.n2580\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__16101\,
            I => \Inst_eia232.Inst_transmitter.n2580\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__16098\,
            I => \Inst_eia232.Inst_transmitter.n2580\
        );

    \I__2061\ : InMux
    port map (
            O => \N__16091\,
            I => \N__16088\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__16088\,
            I => \N__16084\
        );

    \I__2059\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16081\
        );

    \I__2058\ : Span4Mux_s2_h
    port map (
            O => \N__16084\,
            I => \N__16076\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__16081\,
            I => \N__16076\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__16076\,
            I => \N__16073\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__16073\,
            I => \Inst_eia232.Inst_transmitter.n8527\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__16070\,
            I => \N__16065\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__16069\,
            I => \N__16062\
        );

    \I__2052\ : InMux
    port map (
            O => \N__16068\,
            I => \N__16059\
        );

    \I__2051\ : InMux
    port map (
            O => \N__16065\,
            I => \N__16056\
        );

    \I__2050\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16053\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__16059\,
            I => \N__16050\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__16056\,
            I => \N__16047\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__16053\,
            I => \N__16044\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__16050\,
            I => \N__16039\
        );

    \I__2045\ : Span4Mux_s3_h
    port map (
            O => \N__16047\,
            I => \N__16039\
        );

    \I__2044\ : Span4Mux_h
    port map (
            O => \N__16044\,
            I => \N__16036\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__16039\,
            I => \Inst_eia232.id\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__16036\,
            I => \Inst_eia232.id\
        );

    \I__2041\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16028\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__2039\ : Span4Mux_v
    port map (
            O => \N__16025\,
            I => \N__16022\
        );

    \I__2038\ : Span4Mux_v
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__16019\,
            I => \Inst_eia232.Inst_transmitter.n971\
        );

    \I__2036\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16007\
        );

    \I__2035\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16007\
        );

    \I__2034\ : InMux
    port map (
            O => \N__16014\,
            I => \N__16000\
        );

    \I__2033\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16000\
        );

    \I__2032\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16000\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__16007\,
            I => \N__15992\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__16000\,
            I => \N__15992\
        );

    \I__2029\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15977\
        );

    \I__2028\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15974\
        );

    \I__2027\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15971\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__15992\,
            I => \N__15968\
        );

    \I__2025\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15952\
        );

    \I__2024\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15952\
        );

    \I__2023\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15952\
        );

    \I__2022\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15952\
        );

    \I__2021\ : InMux
    port map (
            O => \N__15987\,
            I => \N__15952\
        );

    \I__2020\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15952\
        );

    \I__2019\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15952\
        );

    \I__2018\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15948\
        );

    \I__2017\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15939\
        );

    \I__2016\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15939\
        );

    \I__2015\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15939\
        );

    \I__2014\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15939\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__15977\,
            I => \N__15936\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15931\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15931\
        );

    \I__2010\ : Span4Mux_v
    port map (
            O => \N__15968\,
            I => \N__15928\
        );

    \I__2009\ : InMux
    port map (
            O => \N__15967\,
            I => \N__15925\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__15952\,
            I => \N__15922\
        );

    \I__2007\ : InMux
    port map (
            O => \N__15951\,
            I => \N__15919\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__15948\,
            I => state_1
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__15939\,
            I => state_1
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__15936\,
            I => state_1
        );

    \I__2003\ : Odrv12
    port map (
            O => \N__15931\,
            I => state_1
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__15928\,
            I => state_1
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__15925\,
            I => state_1
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__15922\,
            I => state_1
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__15919\,
            I => state_1
        );

    \I__1998\ : SRMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__15899\,
            I => \N__15896\
        );

    \I__1996\ : Span4Mux_v
    port map (
            O => \N__15896\,
            I => \N__15893\
        );

    \I__1995\ : Span4Mux_s0_h
    port map (
            O => \N__15893\,
            I => \N__15890\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__15890\,
            I => \Inst_eia232.Inst_transmitter.n4712\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__1992\ : CascadeBuf
    port map (
            O => \N__15884\,
            I => \N__15881\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__15881\,
            I => \N__15878\
        );

    \I__1990\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15875\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__15875\,
            I => \GENERIC_FIFO_1.n77\
        );

    \I__1988\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15868\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__15871\,
            I => \N__15865\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__15868\,
            I => \N__15861\
        );

    \I__1985\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15856\
        );

    \I__1984\ : InMux
    port map (
            O => \N__15864\,
            I => \N__15856\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__15861\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__15856\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0\
        );

    \I__1981\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15848\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__15848\,
            I => \N__15844\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__15847\,
            I => \N__15841\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__15844\,
            I => \N__15837\
        );

    \I__1977\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15832\
        );

    \I__1976\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15832\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__15837\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__15832\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4\
        );

    \I__1973\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15824\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__15824\,
            I => \N__15821\
        );

    \I__1971\ : Span4Mux_v
    port map (
            O => \N__15821\,
            I => \N__15818\
        );

    \I__1970\ : Span4Mux_s1_h
    port map (
            O => \N__15818\,
            I => \N__15813\
        );

    \I__1969\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15808\
        );

    \I__1968\ : InMux
    port map (
            O => \N__15816\,
            I => \N__15808\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__15813\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__15808\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__15803\,
            I => \N__15800\
        );

    \I__1964\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15797\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__15797\,
            I => \N__15794\
        );

    \I__1962\ : Span12Mux_s7_v
    port map (
            O => \N__15794\,
            I => \N__15790\
        );

    \I__1961\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15787\
        );

    \I__1960\ : Odrv12
    port map (
            O => \N__15790\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__15787\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__1957\ : CascadeBuf
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__1955\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__1953\ : Span4Mux_s3_h
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__15764\,
            I => \GENERIC_FIFO_1.n71\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__1950\ : CascadeBuf
    port map (
            O => \N__15758\,
            I => \N__15755\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__1948\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15749\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__15743\,
            I => \GENERIC_FIFO_1.n70\
        );

    \I__1944\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__15737\,
            I => \N__15733\
        );

    \I__1942\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15730\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__15733\,
            I => \N__15727\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15724\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__15727\,
            I => \GENERIC_FIFO_1.n8779\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__15724\,
            I => \GENERIC_FIFO_1.n8779\
        );

    \I__1937\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15715\
        );

    \I__1936\ : InMux
    port map (
            O => \N__15718\,
            I => \N__15712\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__15715\,
            I => \valueRegister_0\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__15712\,
            I => \valueRegister_0\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__15707\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_cascade_\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__15704\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9114_cascade_\
        );

    \I__1931\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15698\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__15698\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_0\
        );

    \I__1929\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__1927\ : Span4Mux_s3_h
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__15686\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__1924\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__15671\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9108\
        );

    \I__1920\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15664\
        );

    \I__1919\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15661\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__15664\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__15661\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__15656\,
            I => \N__15652\
        );

    \I__1915\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15648\
        );

    \I__1914\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15645\
        );

    \I__1913\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15642\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__15648\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__15645\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__15642\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16\
        );

    \I__1909\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15624\
        );

    \I__1908\ : InMux
    port map (
            O => \N__15634\,
            I => \N__15624\
        );

    \I__1907\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15624\
        );

    \I__1906\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15621\
        );

    \I__1905\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15618\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__15624\,
            I => \N__15613\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__15621\,
            I => \N__15613\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__15618\,
            I => \Inst_eia232.Inst_receiver.n14_adj_1265\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__15613\,
            I => \Inst_eia232.Inst_receiver.n14_adj_1265\
        );

    \I__1900\ : InMux
    port map (
            O => \N__15608\,
            I => \N__15593\
        );

    \I__1899\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15593\
        );

    \I__1898\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15593\
        );

    \I__1897\ : InMux
    port map (
            O => \N__15605\,
            I => \N__15593\
        );

    \I__1896\ : InMux
    port map (
            O => \N__15604\,
            I => \N__15593\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__15593\,
            I => \Inst_eia232.Inst_receiver.n112\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__15590\,
            I => \Inst_eia232.Inst_receiver.n112_cascade_\
        );

    \I__1893\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15583\
        );

    \I__1892\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15580\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__15583\,
            I => \N__15577\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__15580\,
            I => \Inst_eia232.Inst_receiver.n90\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__15577\,
            I => \Inst_eia232.Inst_receiver.n90\
        );

    \I__1888\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15563\
        );

    \I__1887\ : InMux
    port map (
            O => \N__15571\,
            I => \N__15563\
        );

    \I__1886\ : InMux
    port map (
            O => \N__15570\,
            I => \N__15563\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__15563\,
            I => \N__15559\
        );

    \I__1884\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15556\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__15559\,
            I => \Inst_eia232.Inst_receiver.n5498\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__15556\,
            I => \Inst_eia232.Inst_receiver.n5498\
        );

    \I__1881\ : InMux
    port map (
            O => \N__15551\,
            I => \N__15546\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__15550\,
            I => \N__15542\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__15549\,
            I => \N__15539\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__15546\,
            I => \N__15534\
        );

    \I__1877\ : InMux
    port map (
            O => \N__15545\,
            I => \N__15523\
        );

    \I__1876\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15523\
        );

    \I__1875\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15523\
        );

    \I__1874\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15523\
        );

    \I__1873\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15523\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__15534\,
            I => cmd_6
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__15523\,
            I => cmd_6
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__15518\,
            I => \n5698_cascade_\
        );

    \I__1869\ : InMux
    port map (
            O => \N__15515\,
            I => \N__15512\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__15512\,
            I => \N__15503\
        );

    \I__1867\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15500\
        );

    \I__1866\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15489\
        );

    \I__1865\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15489\
        );

    \I__1864\ : InMux
    port map (
            O => \N__15508\,
            I => \N__15489\
        );

    \I__1863\ : InMux
    port map (
            O => \N__15507\,
            I => \N__15489\
        );

    \I__1862\ : InMux
    port map (
            O => \N__15506\,
            I => \N__15489\
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__15503\,
            I => \nstate_2_N_241_0\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__15500\,
            I => \nstate_2_N_241_0\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__15489\,
            I => \nstate_2_N_241_0\
        );

    \I__1858\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__1856\ : Span4Mux_h
    port map (
            O => \N__15476\,
            I => \N__15472\
        );

    \I__1855\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15469\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__15472\,
            I => \Inst_eia232.xon\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__15469\,
            I => \Inst_eia232.xon\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__15464\,
            I => \Inst_eia232.Inst_receiver.n75_cascade_\
        );

    \I__1851\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__15458\,
            I => \Inst_eia232.Inst_receiver.n5597\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__15455\,
            I => \Inst_eia232.Inst_receiver.n5597_cascade_\
        );

    \I__1848\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__15449\,
            I => \Inst_eia232.xoff\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__15446\,
            I => \Inst_eia232.Inst_receiver.n90_cascade_\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__15443\,
            I => \Inst_eia232.Inst_receiver.n8831_cascade_\
        );

    \I__1844\ : CEMux
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__15437\,
            I => \N__15434\
        );

    \I__1842\ : Span4Mux_h
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__15431\,
            I => \Inst_eia232.Inst_transmitter.n3552\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__15428\,
            I => \Inst_eia232.Inst_receiver.n7_adj_1264_cascade_\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__15425\,
            I => \Inst_eia232.Inst_receiver.n8769_cascade_\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__15422\,
            I => \Inst_eia232.Inst_receiver.n6736_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15416\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__15416\,
            I => \Inst_eia232.Inst_receiver.n8772\
        );

    \I__1835\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15401\
        );

    \I__1834\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15401\
        );

    \I__1833\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15401\
        );

    \I__1832\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15401\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__15401\,
            I => \Inst_eia232.Inst_receiver.bytecount_2\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__15398\,
            I => \N__15392\
        );

    \I__1829\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15388\
        );

    \I__1828\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15379\
        );

    \I__1827\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15379\
        );

    \I__1826\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15379\
        );

    \I__1825\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15379\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__15388\,
            I => \Inst_eia232.Inst_receiver.bytecount_1\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__15379\,
            I => \Inst_eia232.Inst_receiver.bytecount_1\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \Inst_eia232.Inst_receiver.n8582_cascade_\
        );

    \I__1821\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__15368\,
            I => \GENERIC_FIFO_1.n18_adj_1277\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__15365\,
            I => \GENERIC_FIFO_1.n141_cascade_\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__1817\ : CascadeBuf
    port map (
            O => \N__15359\,
            I => \N__15356\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__1815\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__15350\,
            I => \N__15347\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__15344\,
            I => \GENERIC_FIFO_1.n69\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \Inst_eia232.Inst_receiver.n2143_cascade_\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \N__15333\
        );

    \I__1809\ : InMux
    port map (
            O => \N__15337\,
            I => \N__15323\
        );

    \I__1808\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15323\
        );

    \I__1807\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15323\
        );

    \I__1806\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15323\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__15323\,
            I => \Inst_eia232.Inst_receiver.bitcount_1\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__15320\,
            I => \N__15316\
        );

    \I__1803\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15308\
        );

    \I__1802\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15308\
        );

    \I__1801\ : InMux
    port map (
            O => \N__15315\,
            I => \N__15308\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__15308\,
            I => \Inst_eia232.Inst_receiver.bitcount_2\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__15305\,
            I => \N__15301\
        );

    \I__1798\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15296\
        );

    \I__1797\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15296\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__15296\,
            I => \Inst_eia232.Inst_receiver.bitcount_3\
        );

    \I__1795\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15278\
        );

    \I__1794\ : InMux
    port map (
            O => \N__15292\,
            I => \N__15278\
        );

    \I__1793\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15278\
        );

    \I__1792\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15278\
        );

    \I__1791\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15278\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__15278\,
            I => \Inst_eia232.Inst_receiver.bitcount_0\
        );

    \I__1789\ : InMux
    port map (
            O => \N__15275\,
            I => \N__15272\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__15272\,
            I => \GENERIC_FIFO_1.n8650\
        );

    \I__1787\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15266\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__15266\,
            I => \N__15263\
        );

    \I__1785\ : Span4Mux_s2_h
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__15260\,
            I => \GENERIC_FIFO_1.n8681\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \N__15254\
        );

    \I__1782\ : CascadeBuf
    port map (
            O => \N__15254\,
            I => \N__15251\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__15251\,
            I => \N__15248\
        );

    \I__1780\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15245\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__15242\,
            I => \GENERIC_FIFO_1.n78\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__1776\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__15233\,
            I => \GENERIC_FIFO_1.level_9__N_900\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__1773\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15224\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__15221\,
            I => \GENERIC_FIFO_1.n8654\
        );

    \I__1770\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15215\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__15215\,
            I => \GENERIC_FIFO_1.n1418\
        );

    \I__1768\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15209\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__15209\,
            I => \N__15206\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__15206\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_6\
        );

    \I__1765\ : InMux
    port map (
            O => \N__15203\,
            I => \N__15200\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__15200\,
            I => \N__15196\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15193\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__15196\,
            I => \GENERIC_FIFO_1.level_9_N_876_2\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15193\,
            I => \GENERIC_FIFO_1.level_9_N_876_2\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__15188\,
            I => \N__15184\
        );

    \I__1759\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15181\
        );

    \I__1758\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15178\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__15181\,
            I => \N__15175\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__15178\,
            I => \GENERIC_FIFO_1.level_9_N_876_6\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__15175\,
            I => \GENERIC_FIFO_1.level_9_N_876_6\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__1753\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15164\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__15164\,
            I => \N__15160\
        );

    \I__1751\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15157\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__15160\,
            I => \GENERIC_FIFO_1.level_9_N_876_0\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__15157\,
            I => \GENERIC_FIFO_1.level_9_N_876_0\
        );

    \I__1748\ : InMux
    port map (
            O => \N__15152\,
            I => \N__15148\
        );

    \I__1747\ : InMux
    port map (
            O => \N__15151\,
            I => \N__15145\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__15148\,
            I => \GENERIC_FIFO_1.level_9_N_876_8\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__15145\,
            I => \GENERIC_FIFO_1.level_9_N_876_8\
        );

    \I__1744\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15137\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__15137\,
            I => \N__15133\
        );

    \I__1742\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15130\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__15133\,
            I => \GENERIC_FIFO_1.level_9_N_876_5\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__15130\,
            I => \GENERIC_FIFO_1.level_9_N_876_5\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__15125\,
            I => \GENERIC_FIFO_1.n16_adj_1276_cascade_\
        );

    \I__1738\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15118\
        );

    \I__1737\ : InMux
    port map (
            O => \N__15121\,
            I => \N__15115\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__15118\,
            I => \GENERIC_FIFO_1.level_9_N_876_9\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__15115\,
            I => \GENERIC_FIFO_1.level_9_N_876_9\
        );

    \I__1734\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15107\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__15107\,
            I => \GENERIC_FIFO_1.n17_adj_1278\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__1731\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15098\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__15098\,
            I => \N__15095\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__15095\,
            I => \GENERIC_FIFO_1.n1396\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__15092\,
            I => \N__15089\
        );

    \I__1727\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15086\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__15086\,
            I => \GENERIC_FIFO_1.n22\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15083\,
            I => \GENERIC_FIFO_1.n7810\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__1723\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__15074\,
            I => \GENERIC_FIFO_1.n21\
        );

    \I__1721\ : InMux
    port map (
            O => \N__15071\,
            I => \GENERIC_FIFO_1.n7811\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__1719\ : InMux
    port map (
            O => \N__15065\,
            I => \N__15062\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__15062\,
            I => \GENERIC_FIFO_1.n20\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15059\,
            I => \GENERIC_FIFO_1.n7812\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__15056\,
            I => \N__15053\
        );

    \I__1715\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15050\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__15050\,
            I => \GENERIC_FIFO_1.n19\
        );

    \I__1713\ : InMux
    port map (
            O => \N__15047\,
            I => \GENERIC_FIFO_1.n7813\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__15044\,
            I => \N__15041\
        );

    \I__1711\ : InMux
    port map (
            O => \N__15041\,
            I => \N__15038\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__15038\,
            I => \N__15035\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__15035\,
            I => \GENERIC_FIFO_1.n18_adj_1275\
        );

    \I__1708\ : InMux
    port map (
            O => \N__15032\,
            I => \GENERIC_FIFO_1.n7814\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__15029\,
            I => \N__15026\
        );

    \I__1706\ : InMux
    port map (
            O => \N__15026\,
            I => \N__15023\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__15023\,
            I => \GENERIC_FIFO_1.n17\
        );

    \I__1704\ : InMux
    port map (
            O => \N__15020\,
            I => \GENERIC_FIFO_1.n7815\
        );

    \I__1703\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__15014\,
            I => \GENERIC_FIFO_1.n16_adj_1273\
        );

    \I__1701\ : InMux
    port map (
            O => \N__15011\,
            I => \bfn_2_14_0_\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15008\,
            I => \GENERIC_FIFO_1.n7817\
        );

    \I__1699\ : InMux
    port map (
            O => \N__15005\,
            I => \N__15002\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__15002\,
            I => \GENERIC_FIFO_1.n15\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__14999\,
            I => \GENERIC_FIFO_1.n18_cascade_\
        );

    \I__1696\ : CEMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__14993\,
            I => \N__14988\
        );

    \I__1694\ : SRMux
    port map (
            O => \N__14992\,
            I => \N__14985\
        );

    \I__1693\ : SRMux
    port map (
            O => \N__14991\,
            I => \N__14982\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__14988\,
            I => \N__14978\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__14985\,
            I => \N__14975\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__14982\,
            I => \N__14972\
        );

    \I__1689\ : CEMux
    port map (
            O => \N__14981\,
            I => \N__14968\
        );

    \I__1688\ : Span4Mux_s1_h
    port map (
            O => \N__14978\,
            I => \N__14963\
        );

    \I__1687\ : Span4Mux_h
    port map (
            O => \N__14975\,
            I => \N__14963\
        );

    \I__1686\ : Span4Mux_h
    port map (
            O => \N__14972\,
            I => \N__14960\
        );

    \I__1685\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14957\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__14968\,
            I => \GENERIC_FIFO_1.fifo_memory_N_983\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__14963\,
            I => \GENERIC_FIFO_1.fifo_memory_N_983\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__14960\,
            I => \GENERIC_FIFO_1.fifo_memory_N_983\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__14957\,
            I => \GENERIC_FIFO_1.fifo_memory_N_983\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__14948\,
            I => \N__14945\
        );

    \I__1679\ : CascadeBuf
    port map (
            O => \N__14945\,
            I => \N__14942\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__14942\,
            I => \N__14939\
        );

    \I__1677\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14935\
        );

    \I__1676\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14931\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__14935\,
            I => \N__14926\
        );

    \I__1674\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14923\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__14931\,
            I => \N__14920\
        );

    \I__1672\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14915\
        );

    \I__1671\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14915\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__14926\,
            I => \N__14912\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__14923\,
            I => \GENERIC_FIFO_1.write_pointer_4\
        );

    \I__1668\ : Odrv12
    port map (
            O => \N__14920\,
            I => \GENERIC_FIFO_1.write_pointer_4\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__14915\,
            I => \GENERIC_FIFO_1.write_pointer_4\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__14912\,
            I => \GENERIC_FIFO_1.write_pointer_4\
        );

    \I__1665\ : InMux
    port map (
            O => \N__14903\,
            I => \N__14900\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__14900\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_4\
        );

    \I__1663\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14894\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__14891\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_5\
        );

    \I__1660\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__1658\ : Odrv12
    port map (
            O => \N__14882\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n11\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__1656\ : CascadeBuf
    port map (
            O => \N__14876\,
            I => \N__14872\
        );

    \I__1655\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14869\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__14872\,
            I => \N__14865\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__14869\,
            I => \N__14860\
        );

    \I__1652\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14857\
        );

    \I__1651\ : InMux
    port map (
            O => \N__14865\,
            I => \N__14854\
        );

    \I__1650\ : InMux
    port map (
            O => \N__14864\,
            I => \N__14851\
        );

    \I__1649\ : InMux
    port map (
            O => \N__14863\,
            I => \N__14848\
        );

    \I__1648\ : Span4Mux_s2_v
    port map (
            O => \N__14860\,
            I => \N__14843\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__14857\,
            I => \N__14843\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__14854\,
            I => \N__14840\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__14851\,
            I => \GENERIC_FIFO_1.write_pointer_5\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__14848\,
            I => \GENERIC_FIFO_1.write_pointer_5\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__14843\,
            I => \GENERIC_FIFO_1.write_pointer_5\
        );

    \I__1642\ : Odrv12
    port map (
            O => \N__14840\,
            I => \GENERIC_FIFO_1.write_pointer_5\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__14831\,
            I => \GENERIC_FIFO_1.n16_cascade_\
        );

    \I__1640\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__14825\,
            I => \GENERIC_FIFO_1.n20_adj_1274\
        );

    \I__1638\ : SRMux
    port map (
            O => \N__14822\,
            I => \N__14818\
        );

    \I__1637\ : SRMux
    port map (
            O => \N__14821\,
            I => \N__14815\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__14818\,
            I => \GENERIC_FIFO_1.n4721\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__14815\,
            I => \GENERIC_FIFO_1.n4721\
        );

    \I__1634\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__14807\,
            I => \N__14804\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__14804\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105\
        );

    \I__1631\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__14798\,
            I => \N__14795\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__14795\,
            I => \GENERIC_FIFO_1.level_9_N_925_0\
        );

    \I__1628\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14789\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__14789\,
            I => \GENERIC_FIFO_1.n24\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__1625\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__14780\,
            I => \GENERIC_FIFO_1.n23\
        );

    \I__1623\ : InMux
    port map (
            O => \N__14777\,
            I => \GENERIC_FIFO_1.n7809\
        );

    \I__1622\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14770\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14773\,
            I => \N__14767\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__14770\,
            I => \N__14764\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__14767\,
            I => \maskRegister_5\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__14764\,
            I => \maskRegister_5\
        );

    \I__1617\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14755\
        );

    \I__1616\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14746\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__14755\,
            I => \N__14743\
        );

    \I__1614\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14738\
        );

    \I__1613\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14738\
        );

    \I__1612\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14729\
        );

    \I__1611\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14729\
        );

    \I__1610\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14729\
        );

    \I__1609\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14729\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14724\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__14743\,
            I => \N__14724\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__14738\,
            I => \Inst_eia232.Inst_transmitter.n6703\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__14729\,
            I => \Inst_eia232.Inst_transmitter.n6703\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__14724\,
            I => \Inst_eia232.Inst_transmitter.n6703\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__14717\,
            I => \N__14714\
        );

    \I__1602\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__14711\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_5\
        );

    \I__1600\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__14705\,
            I => \N__14702\
        );

    \I__1598\ : Span4Mux_v
    port map (
            O => \N__14702\,
            I => \N__14698\
        );

    \I__1597\ : InMux
    port map (
            O => \N__14701\,
            I => \N__14695\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__14698\,
            I => \Inst_eia232.Inst_transmitter.byte_5\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__14695\,
            I => \Inst_eia232.Inst_transmitter.byte_5\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__14690\,
            I => \GENERIC_FIFO_1.n8677_cascade_\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__14687\,
            I => \GENERIC_FIFO_1.n1396_cascade_\
        );

    \I__1592\ : SRMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__14681\,
            I => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4743\
        );

    \I__1590\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14675\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__14675\,
            I => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_0\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__1587\ : CascadeBuf
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__1585\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14658\
        );

    \I__1584\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14651\
        );

    \I__1583\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14651\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__14658\,
            I => \N__14648\
        );

    \I__1581\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14645\
        );

    \I__1580\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14642\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__14651\,
            I => \N__14639\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__14648\,
            I => \N__14636\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__14645\,
            I => \GENERIC_FIFO_1.write_pointer_8\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14642\,
            I => \GENERIC_FIFO_1.write_pointer_8\
        );

    \I__1575\ : Odrv12
    port map (
            O => \N__14639\,
            I => \GENERIC_FIFO_1.write_pointer_8\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__14636\,
            I => \GENERIC_FIFO_1.write_pointer_8\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__1572\ : CascadeBuf
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__1570\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14612\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__14617\,
            I => \N__14608\
        );

    \I__1568\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14603\
        );

    \I__1567\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14603\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__14612\,
            I => \N__14600\
        );

    \I__1565\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14597\
        );

    \I__1564\ : InMux
    port map (
            O => \N__14608\,
            I => \N__14594\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__14603\,
            I => \N__14591\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__14600\,
            I => \N__14588\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__14597\,
            I => \GENERIC_FIFO_1.write_pointer_9\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__14594\,
            I => \GENERIC_FIFO_1.write_pointer_9\
        );

    \I__1559\ : Odrv12
    port map (
            O => \N__14591\,
            I => \GENERIC_FIFO_1.write_pointer_9\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__14588\,
            I => \GENERIC_FIFO_1.write_pointer_9\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__14579\,
            I => \N__14576\
        );

    \I__1556\ : CascadeBuf
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__14573\,
            I => \N__14568\
        );

    \I__1554\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14563\
        );

    \I__1553\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14560\
        );

    \I__1552\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14557\
        );

    \I__1551\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14554\
        );

    \I__1550\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14551\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__14563\,
            I => \N__14546\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__14560\,
            I => \N__14546\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__14557\,
            I => \N__14543\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__14554\,
            I => \GENERIC_FIFO_1.write_pointer_7\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__14551\,
            I => \GENERIC_FIFO_1.write_pointer_7\
        );

    \I__1544\ : Odrv12
    port map (
            O => \N__14546\,
            I => \GENERIC_FIFO_1.write_pointer_7\
        );

    \I__1543\ : Odrv12
    port map (
            O => \N__14543\,
            I => \GENERIC_FIFO_1.write_pointer_7\
        );

    \I__1542\ : InMux
    port map (
            O => \N__14534\,
            I => \GENERIC_FIFO_1.n7930\
        );

    \I__1541\ : InMux
    port map (
            O => \N__14531\,
            I => \GENERIC_FIFO_1.n7931\
        );

    \I__1540\ : InMux
    port map (
            O => \N__14528\,
            I => \GENERIC_FIFO_1.n7932\
        );

    \I__1539\ : InMux
    port map (
            O => \N__14525\,
            I => \GENERIC_FIFO_1.n7933\
        );

    \I__1538\ : InMux
    port map (
            O => \N__14522\,
            I => \GENERIC_FIFO_1.n7934\
        );

    \I__1537\ : InMux
    port map (
            O => \N__14519\,
            I => \GENERIC_FIFO_1.n7935\
        );

    \I__1536\ : InMux
    port map (
            O => \N__14516\,
            I => \bfn_2_9_0_\
        );

    \I__1535\ : InMux
    port map (
            O => \N__14513\,
            I => \GENERIC_FIFO_1.n7937\
        );

    \I__1534\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14504\
        );

    \I__1533\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14504\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__14504\,
            I => \disabledGroupsReg_3\
        );

    \I__1531\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14497\
        );

    \I__1530\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14494\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__14497\,
            I => \N__14491\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__14494\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_2\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__14491\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_2\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__14486\,
            I => \N__14483\
        );

    \I__1525\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14477\
        );

    \I__1524\ : InMux
    port map (
            O => \N__14482\,
            I => \N__14477\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__14477\,
            I => \disabledGroupsReg_2\
        );

    \I__1522\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14471\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__14471\,
            I => \N__14468\
        );

    \I__1520\ : Span4Mux_s2_h
    port map (
            O => \N__14468\,
            I => \N__14464\
        );

    \I__1519\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14461\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__14464\,
            I => \Inst_eia232.Inst_transmitter.byte_7\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__14461\,
            I => \Inst_eia232.Inst_transmitter.byte_7\
        );

    \I__1516\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__14450\,
            I => \N__14447\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__14447\,
            I => outputdata_7
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__14444\,
            I => \N__14440\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__14443\,
            I => \N__14437\
        );

    \I__1510\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14432\
        );

    \I__1509\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14432\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__14432\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_7\
        );

    \I__1507\ : InMux
    port map (
            O => \N__14429\,
            I => \bfn_2_8_0_\
        );

    \I__1506\ : InMux
    port map (
            O => \N__14426\,
            I => \GENERIC_FIFO_1.n7929\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__14423\,
            I => \N__14419\
        );

    \I__1504\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14405\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14405\
        );

    \I__1502\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14405\
        );

    \I__1501\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14400\
        );

    \I__1500\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14400\
        );

    \I__1499\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14391\
        );

    \I__1498\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14391\
        );

    \I__1497\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14391\
        );

    \I__1496\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14391\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__14405\,
            I => bytes_0
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__14400\,
            I => bytes_0
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__14391\,
            I => bytes_0
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__14384\,
            I => \Inst_eia232.Inst_transmitter.n3652_cascade_\
        );

    \I__1491\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14378\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__14378\,
            I => n1336
        );

    \I__1489\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14372\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__14372\,
            I => \N__14369\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__14369\,
            I => \N__14366\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__14366\,
            I => outputdata_1
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__14363\,
            I => \N__14359\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14362\,
            I => \N__14356\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14353\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14350\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__14353\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_1\
        );

    \I__1480\ : Odrv12
    port map (
            O => \N__14350\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_1\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14342\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14339\
        );

    \I__1477\ : Sp12to4
    port map (
            O => \N__14339\,
            I => \N__14336\
        );

    \I__1476\ : Odrv12
    port map (
            O => \N__14336\,
            I => outputdata_2
        );

    \I__1475\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14329\
        );

    \I__1474\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14326\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__14329\,
            I => \N__14323\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__14326\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_2\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__14323\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_2\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__14318\,
            I => \N__14315\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14312\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__14312\,
            I => \N__14309\
        );

    \I__1467\ : Span12Mux_s11_v
    port map (
            O => \N__14309\,
            I => \N__14306\
        );

    \I__1466\ : Odrv12
    port map (
            O => \N__14306\,
            I => outputdata_3
        );

    \I__1465\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14299\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14296\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__14299\,
            I => \N__14293\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__14296\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_3\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__14293\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_3\
        );

    \I__1460\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14285\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__14285\,
            I => \N__14282\
        );

    \I__1458\ : Span4Mux_s2_h
    port map (
            O => \N__14282\,
            I => \N__14279\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__14279\,
            I => outputdata_6
        );

    \I__1456\ : InMux
    port map (
            O => \N__14276\,
            I => \N__14272\
        );

    \I__1455\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14269\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__14272\,
            I => \N__14266\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__14269\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_6\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__14266\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_6\
        );

    \I__1451\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14257\
        );

    \I__1450\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14254\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__14257\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_1\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__14254\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_1\
        );

    \I__1447\ : InMux
    port map (
            O => \N__14249\,
            I => \N__14243\
        );

    \I__1446\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14243\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__14243\,
            I => \disabledGroupsReg_1\
        );

    \I__1444\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14236\
        );

    \I__1443\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14233\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__14236\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_3\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__14233\,
            I => \Inst_eia232.Inst_transmitter.disabledBuffer_3\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__14228\,
            I => \n1320_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14221\
        );

    \I__1438\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14218\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__14221\,
            I => \dataBuffer_28\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__14218\,
            I => \dataBuffer_28\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__14213\,
            I => \Inst_eia232.Inst_transmitter.n8756_cascade_\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14207\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__14204\,
            I => \N__14201\
        );

    \I__1431\ : Span4Mux_h
    port map (
            O => \N__14201\,
            I => \N__14198\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__14198\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_4\
        );

    \I__1429\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__14192\,
            I => \Inst_eia232.Inst_transmitter.byte_4\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__14189\,
            I => \state_1_N_371_1_cascade_\
        );

    \I__1426\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14183\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__14183\,
            I => \Inst_eia232.Inst_transmitter.n1\
        );

    \I__1424\ : InMux
    port map (
            O => \N__14180\,
            I => \N__14166\
        );

    \I__1423\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14166\
        );

    \I__1422\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14166\
        );

    \I__1421\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14161\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14161\
        );

    \I__1419\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14154\
        );

    \I__1418\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14154\
        );

    \I__1417\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14154\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__14166\,
            I => bytes_1
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__14161\,
            I => bytes_1
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__14154\,
            I => bytes_1
        );

    \I__1413\ : InMux
    port map (
            O => \N__14147\,
            I => \N__14137\
        );

    \I__1412\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14137\
        );

    \I__1411\ : InMux
    port map (
            O => \N__14145\,
            I => \N__14134\
        );

    \I__1410\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14131\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14143\,
            I => \N__14126\
        );

    \I__1408\ : InMux
    port map (
            O => \N__14142\,
            I => \N__14126\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__14137\,
            I => bytes_2
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__14134\,
            I => bytes_2
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__14131\,
            I => bytes_2
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__14126\,
            I => bytes_2
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__14117\,
            I => \Inst_eia232.Inst_transmitter.n9218_cascade_\
        );

    \I__1402\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14111\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__14111\,
            I => \Inst_eia232.Inst_transmitter.n3\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14105\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__14105\,
            I => \N__14102\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__14102\,
            I => disabled
        );

    \I__1397\ : CEMux
    port map (
            O => \N__14099\,
            I => \N__14096\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__14096\,
            I => \N__14093\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__14093\,
            I => \Inst_eia232.Inst_transmitter.n6745\
        );

    \I__1394\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14083\
        );

    \I__1393\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14083\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14080\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__14083\,
            I => \state_1_N_371_1\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14080\,
            I => \state_1_N_371_1\
        );

    \I__1389\ : CEMux
    port map (
            O => \N__14075\,
            I => \N__14072\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__14072\,
            I => \N__14068\
        );

    \I__1387\ : CEMux
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__1386\ : Span4Mux_s3_v
    port map (
            O => \N__14068\,
            I => \N__14060\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__14065\,
            I => \N__14060\
        );

    \I__1384\ : Span4Mux_h
    port map (
            O => \N__14060\,
            I => \N__14056\
        );

    \I__1383\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14053\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__14056\,
            I => \Inst_eia232.Inst_transmitter.n3652\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__14053\,
            I => \Inst_eia232.Inst_transmitter.n3652\
        );

    \I__1380\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14045\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__14045\,
            I => \Inst_eia232.Inst_transmitter.n1323\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__14042\,
            I => \Inst_eia232.Inst_transmitter.n3632_cascade_\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14036\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__14036\,
            I => \Inst_eia232.Inst_transmitter.byte_6\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__14033\,
            I => \N__14029\
        );

    \I__1374\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__1373\ : InMux
    port map (
            O => \N__14029\,
            I => \N__14023\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__14026\,
            I => \dataBuffer_18\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__14023\,
            I => \dataBuffer_18\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__14018\,
            I => \Inst_eia232.Inst_transmitter.n8851_cascade_\
        );

    \I__1369\ : InMux
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__1367\ : Odrv12
    port map (
            O => \N__14009\,
            I => \Inst_eia232.Inst_transmitter.byte_2\
        );

    \I__1366\ : InMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__14003\,
            I => \Inst_eia232.Inst_transmitter.byte_1\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__14000\,
            I => \n4248_cascade_\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__13997\,
            I => \n1336_cascade_\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__13994\,
            I => \N__13991\
        );

    \I__1361\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13987\
        );

    \I__1360\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13984\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__13987\,
            I => \dataBuffer_25\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__13984\,
            I => \dataBuffer_25\
        );

    \I__1357\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13976\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__13976\,
            I => \Inst_eia232.Inst_transmitter.n8847\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__1354\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__13967\,
            I => n4248
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__1351\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13954\
        );

    \I__1350\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13951\
        );

    \I__1349\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13946\
        );

    \I__1348\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13946\
        );

    \I__1347\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13943\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__13954\,
            I => \N__13938\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__13951\,
            I => \N__13938\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__13946\,
            I => n1320
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__13943\,
            I => n1320
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__13938\,
            I => n1320
        );

    \I__1341\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13925\
        );

    \I__1340\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13925\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__13925\,
            I => \dataBuffer_22\
        );

    \I__1338\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13916\
        );

    \I__1337\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13916\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__13916\,
            I => \dataBuffer_30\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__13913\,
            I => \N__13909\
        );

    \I__1334\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13906\
        );

    \I__1333\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13903\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__13906\,
            I => \dataBuffer_24\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__13903\,
            I => \dataBuffer_24\
        );

    \I__1330\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__1328\ : Odrv12
    port map (
            O => \N__13892\,
            I => \Inst_eia232.Inst_transmitter.byte_0\
        );

    \I__1327\ : InMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__13883\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_8\
        );

    \I__1324\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__1322\ : Span4Mux_v
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__13871\,
            I => \Inst_eia232.Inst_transmitter.dataBuffer_0\
        );

    \I__1320\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__13865\,
            I => \Inst_eia232.Inst_transmitter.n3571\
        );

    \I__1318\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13858\
        );

    \I__1317\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13855\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__13858\,
            I => \dataBuffer_19\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__13855\,
            I => \dataBuffer_19\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__13850\,
            I => \Inst_eia232.Inst_transmitter.n8854_cascade_\
        );

    \I__1313\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__13844\,
            I => \Inst_eia232.Inst_transmitter.byte_3\
        );

    \I__1311\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13837\
        );

    \I__1310\ : InMux
    port map (
            O => \N__13840\,
            I => \N__13834\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__13837\,
            I => \dataBuffer_14\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__13834\,
            I => \dataBuffer_14\
        );

    \I__1307\ : InMux
    port map (
            O => \N__13829\,
            I => \GENERIC_FIFO_1.n7826\
        );

    \I__1306\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13823\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__13820\,
            I => \GENERIC_FIFO_1.n3\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__13817\,
            I => \n4005_cascade_\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__1301\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13808\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__13808\,
            I => \N__13805\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__13805\,
            I => \GENERIC_FIFO_1.n12\
        );

    \I__1298\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13799\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__13799\,
            I => \N__13796\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__13796\,
            I => \GENERIC_FIFO_1.n11\
        );

    \I__1295\ : InMux
    port map (
            O => \N__13793\,
            I => \GENERIC_FIFO_1.n7818\
        );

    \I__1294\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13787\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__13787\,
            I => \N__13784\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__13784\,
            I => \GENERIC_FIFO_1.n10\
        );

    \I__1291\ : InMux
    port map (
            O => \N__13781\,
            I => \GENERIC_FIFO_1.n7819\
        );

    \I__1290\ : InMux
    port map (
            O => \N__13778\,
            I => \N__13775\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__13775\,
            I => \N__13772\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__13772\,
            I => \GENERIC_FIFO_1.n9\
        );

    \I__1287\ : InMux
    port map (
            O => \N__13769\,
            I => \GENERIC_FIFO_1.n7820\
        );

    \I__1286\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13763\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__13763\,
            I => \N__13760\
        );

    \I__1284\ : Span4Mux_s1_h
    port map (
            O => \N__13760\,
            I => \N__13757\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__13757\,
            I => \GENERIC_FIFO_1.n8\
        );

    \I__1282\ : InMux
    port map (
            O => \N__13754\,
            I => \GENERIC_FIFO_1.n7821\
        );

    \I__1281\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13748\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__13748\,
            I => \N__13745\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__13745\,
            I => \GENERIC_FIFO_1.n7\
        );

    \I__1278\ : InMux
    port map (
            O => \N__13742\,
            I => \GENERIC_FIFO_1.n7822\
        );

    \I__1277\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__13736\,
            I => \N__13733\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__13733\,
            I => \GENERIC_FIFO_1.n6\
        );

    \I__1274\ : InMux
    port map (
            O => \N__13730\,
            I => \GENERIC_FIFO_1.n7823\
        );

    \I__1273\ : InMux
    port map (
            O => \N__13727\,
            I => \N__13724\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__13724\,
            I => \N__13721\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__13721\,
            I => \GENERIC_FIFO_1.n5\
        );

    \I__1270\ : InMux
    port map (
            O => \N__13718\,
            I => \GENERIC_FIFO_1.n7824\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__13715\,
            I => \N__13712\
        );

    \I__1268\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13709\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__13706\,
            I => \GENERIC_FIFO_1.n4\
        );

    \I__1265\ : InMux
    port map (
            O => \N__13703\,
            I => \bfn_1_16_0_\
        );

    \I__1264\ : InMux
    port map (
            O => \N__13700\,
            I => \GENERIC_FIFO_1.n7830\
        );

    \I__1263\ : InMux
    port map (
            O => \N__13697\,
            I => \GENERIC_FIFO_1.n7831\
        );

    \I__1262\ : InMux
    port map (
            O => \N__13694\,
            I => \GENERIC_FIFO_1.n7832\
        );

    \I__1261\ : InMux
    port map (
            O => \N__13691\,
            I => \GENERIC_FIFO_1.n7833\
        );

    \I__1260\ : InMux
    port map (
            O => \N__13688\,
            I => \bfn_1_14_0_\
        );

    \I__1259\ : InMux
    port map (
            O => \N__13685\,
            I => \GENERIC_FIFO_1.n7835\
        );

    \I__1258\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13678\
        );

    \I__1257\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13675\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__13678\,
            I => \N__13672\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__13675\,
            I => \GENERIC_FIFO_1.level_9_N_876_7\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__13672\,
            I => \GENERIC_FIFO_1.level_9_N_876_7\
        );

    \I__1253\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13663\
        );

    \I__1252\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13660\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__13663\,
            I => \GENERIC_FIFO_1.level_9_N_876_1\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__13660\,
            I => \GENERIC_FIFO_1.level_9_N_876_1\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__13655\,
            I => \N__13651\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__13654\,
            I => \N__13648\
        );

    \I__1247\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13645\
        );

    \I__1246\ : InMux
    port map (
            O => \N__13648\,
            I => \N__13642\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__13645\,
            I => \GENERIC_FIFO_1.level_9_N_876_4\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__13642\,
            I => \GENERIC_FIFO_1.level_9_N_876_4\
        );

    \I__1243\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13633\
        );

    \I__1242\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13630\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__13633\,
            I => \GENERIC_FIFO_1.level_9_N_876_3\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__13630\,
            I => \GENERIC_FIFO_1.level_9_N_876_3\
        );

    \I__1239\ : InMux
    port map (
            O => \N__13625\,
            I => \GENERIC_FIFO_1.n7840\
        );

    \I__1238\ : InMux
    port map (
            O => \N__13622\,
            I => \GENERIC_FIFO_1.n7841\
        );

    \I__1237\ : InMux
    port map (
            O => \N__13619\,
            I => \GENERIC_FIFO_1.n7842\
        );

    \I__1236\ : InMux
    port map (
            O => \N__13616\,
            I => \bfn_1_12_0_\
        );

    \I__1235\ : InMux
    port map (
            O => \N__13613\,
            I => \GENERIC_FIFO_1.n7844\
        );

    \I__1234\ : InMux
    port map (
            O => \N__13610\,
            I => \GENERIC_FIFO_1.n7827\
        );

    \I__1233\ : InMux
    port map (
            O => \N__13607\,
            I => \GENERIC_FIFO_1.n7828\
        );

    \I__1232\ : InMux
    port map (
            O => \N__13604\,
            I => \GENERIC_FIFO_1.n7829\
        );

    \I__1231\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13598\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__13598\,
            I => \N__13595\
        );

    \I__1229\ : Span4Mux_s3_h
    port map (
            O => \N__13595\,
            I => \N__13592\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__13592\,
            I => outputdata_0
        );

    \I__1227\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__13586\,
            I => \N__13583\
        );

    \I__1225\ : Odrv12
    port map (
            O => \N__13583\,
            I => outputdata_4
        );

    \I__1224\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13577\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__13577\,
            I => \N__13574\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__13574\,
            I => outputdata_5
        );

    \I__1221\ : InMux
    port map (
            O => \N__13571\,
            I => \N__13568\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__13568\,
            I => \N__13565\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__13562\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_1\
        );

    \I__1217\ : IoInMux
    port map (
            O => \N__13559\,
            I => \N__13556\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__13556\,
            I => \N__13553\
        );

    \I__1215\ : Span4Mux_s0_h
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__13550\,
            I => tx_c
        );

    \I__1213\ : InMux
    port map (
            O => \N__13547\,
            I => \bfn_1_11_0_\
        );

    \I__1212\ : InMux
    port map (
            O => \N__13544\,
            I => \GENERIC_FIFO_1.n7836\
        );

    \I__1211\ : InMux
    port map (
            O => \N__13541\,
            I => \GENERIC_FIFO_1.n7837\
        );

    \I__1210\ : InMux
    port map (
            O => \N__13538\,
            I => \GENERIC_FIFO_1.n7838\
        );

    \I__1209\ : InMux
    port map (
            O => \N__13535\,
            I => \GENERIC_FIFO_1.n7839\
        );

    \I__1208\ : InMux
    port map (
            O => \N__13532\,
            I => \N__13525\
        );

    \I__1207\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13525\
        );

    \I__1206\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13522\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__13525\,
            I => \Inst_eia232.Inst_transmitter.counter_3\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__13522\,
            I => \Inst_eia232.Inst_transmitter.counter_3\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__13517\,
            I => \Inst_eia232.Inst_transmitter.n2201_cascade_\
        );

    \I__1202\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13508\
        );

    \I__1201\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13508\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__13508\,
            I => \Inst_eia232.Inst_transmitter.counter_4\
        );

    \I__1199\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13502\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__13502\,
            I => \Inst_eia232.Inst_transmitter.n8642\
        );

    \I__1197\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13484\
        );

    \I__1196\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13484\
        );

    \I__1195\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13484\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13484\
        );

    \I__1193\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13484\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__13484\,
            I => \Inst_eia232.Inst_transmitter.counter_1\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__13481\,
            I => \N__13476\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__13480\,
            I => \N__13472\
        );

    \I__1189\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13465\
        );

    \I__1188\ : InMux
    port map (
            O => \N__13476\,
            I => \N__13465\
        );

    \I__1187\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13465\
        );

    \I__1186\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13462\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__13465\,
            I => \Inst_eia232.Inst_transmitter.counter_2\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__13462\,
            I => \Inst_eia232.Inst_transmitter.counter_2\
        );

    \I__1183\ : CEMux
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__1181\ : Span4Mux_v
    port map (
            O => \N__13451\,
            I => \N__13448\
        );

    \I__1180\ : Span4Mux_s0_h
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__13445\,
            I => \Inst_eia232.Inst_transmitter.n3594\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__13442\,
            I => \Inst_eia232.Inst_transmitter.n3594_cascade_\
        );

    \I__1177\ : SRMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__1175\ : Span4Mux_s1_h
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__13430\,
            I => \Inst_eia232.Inst_transmitter.n4719\
        );

    \I__1173\ : CEMux
    port map (
            O => \N__13427\,
            I => \N__13423\
        );

    \I__1172\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13420\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__13423\,
            I => \N__13415\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__13420\,
            I => \N__13415\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__13415\,
            I => n3615
        );

    \I__1168\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13404\
        );

    \I__1167\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13401\
        );

    \I__1166\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13392\
        );

    \I__1165\ : InMux
    port map (
            O => \N__13409\,
            I => \N__13392\
        );

    \I__1164\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13392\
        );

    \I__1163\ : InMux
    port map (
            O => \N__13407\,
            I => \N__13392\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__13404\,
            I => \N__13389\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__13401\,
            I => \Inst_eia232.Inst_transmitter.counter_0\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__13392\,
            I => \Inst_eia232.Inst_transmitter.counter_0\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__13389\,
            I => \Inst_eia232.Inst_transmitter.counter_0\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__13382\,
            I => \n9_cascade_\
        );

    \I__1157\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13373\
        );

    \I__1156\ : InMux
    port map (
            O => \N__13378\,
            I => \N__13373\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__13373\,
            I => \Inst_eia232.Inst_transmitter.bits_3\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__13370\,
            I => \N__13366\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__13369\,
            I => \N__13362\
        );

    \I__1152\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13355\
        );

    \I__1151\ : InMux
    port map (
            O => \N__13365\,
            I => \N__13355\
        );

    \I__1150\ : InMux
    port map (
            O => \N__13362\,
            I => \N__13355\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__13355\,
            I => \Inst_eia232.Inst_transmitter.bits_2\
        );

    \I__1148\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13349\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__13349\,
            I => n3493
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__13346\,
            I => \n3493_cascade_\
        );

    \I__1145\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13340\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__13340\,
            I => \N__13337\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__13337\,
            I => n6749
        );

    \I__1142\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13327\
        );

    \I__1141\ : InMux
    port map (
            O => \N__13333\,
            I => \N__13320\
        );

    \I__1140\ : InMux
    port map (
            O => \N__13332\,
            I => \N__13320\
        );

    \I__1139\ : InMux
    port map (
            O => \N__13331\,
            I => \N__13320\
        );

    \I__1138\ : InMux
    port map (
            O => \N__13330\,
            I => \N__13317\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__13327\,
            I => \N__13312\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__13320\,
            I => \N__13312\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__13317\,
            I => \Inst_eia232.Inst_transmitter.bits_0\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__13312\,
            I => \Inst_eia232.Inst_transmitter.bits_0\
        );

    \I__1133\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13295\
        );

    \I__1132\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13295\
        );

    \I__1131\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13295\
        );

    \I__1130\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13295\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__13295\,
            I => \Inst_eia232.Inst_transmitter.bits_1\
        );

    \I__1128\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13288\
        );

    \I__1127\ : CEMux
    port map (
            O => \N__13291\,
            I => \N__13285\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__13288\,
            I => \N__13282\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__13285\,
            I => n4082
        );

    \I__1124\ : Odrv12
    port map (
            O => \N__13282\,
            I => n4082
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__13277\,
            I => \n234_cascade_\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__13274\,
            I => \N__13270\
        );

    \I__1121\ : InMux
    port map (
            O => \N__13273\,
            I => \N__13267\
        );

    \I__1120\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13264\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__13267\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_9\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__13264\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_9\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__13259\,
            I => \N__13256\
        );

    \I__1116\ : InMux
    port map (
            O => \N__13256\,
            I => \N__13253\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__13253\,
            I => n234
        );

    \I__1114\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13244\
        );

    \I__1113\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13244\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__13244\,
            I => \byteDone\
        );

    \I__1111\ : InMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__13238\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_6\
        );

    \I__1109\ : InMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__13232\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_5\
        );

    \I__1107\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__13226\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_4\
        );

    \I__1105\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__13220\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_3\
        );

    \I__1103\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__13214\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_2\
        );

    \I__1101\ : InMux
    port map (
            O => \N__13211\,
            I => \N__13208\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__13208\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_7\
        );

    \I__1099\ : InMux
    port map (
            O => \N__13205\,
            I => \N__13202\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__13202\,
            I => \Inst_eia232.Inst_transmitter.txBuffer_8\
        );

    \INVInst_core.Inst_sync.synchronizedInput180_i0C\ : INV
    port map (
            O => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            I => \N__37605\
        );

    \INVInst_core.Inst_sync.synchronizedInput180_i4C\ : INV
    port map (
            O => \INVInst_core.Inst_sync.synchronizedInput180_i4C_net\,
            I => \N__37594\
        );

    \IN_MUX_bfv_6_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_1_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7921\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7906\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7891\,
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7876\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_sampler.n7955\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_sampler.n7963\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_controller.n7852\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Inst_core.Inst_controller.n7860\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \GENERIC_FIFO_1.n7843\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \GENERIC_FIFO_1.n7936\,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \GENERIC_FIFO_1.n7816\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \GENERIC_FIFO_1.n7825\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \GENERIC_FIFO_1.n7944_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \GENERIC_FIFO_1.n7834\,
            carryinitout => \bfn_1_14_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.paused_91_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15482\,
            lcout => \Inst_eia232.Inst_transmitter.paused\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37515\,
            ce => \N__15440\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.bits__i0_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13330\,
            in2 => \_gnd_net_\,
            in3 => \N__13292\,
            lcout => \Inst_eia232.Inst_transmitter.bits_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37506\,
            ce => 'H',
            sr => \N__16822\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i7_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14708\,
            in1 => \N__13211\,
            in2 => \_gnd_net_\,
            in3 => \N__16794\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i6_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16791\,
            in1 => \N__14195\,
            in2 => \_gnd_net_\,
            in3 => \N__13241\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i5_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13847\,
            in1 => \N__13235\,
            in2 => \_gnd_net_\,
            in3 => \N__16793\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i4_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16790\,
            in1 => \N__14015\,
            in2 => \_gnd_net_\,
            in3 => \N__13229\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i3_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16823\,
            in1 => \N__13223\,
            in2 => \_gnd_net_\,
            in3 => \N__14006\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i2_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16789\,
            in1 => \N__13898\,
            in2 => \_gnd_net_\,
            in3 => \N__13217\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i8_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14039\,
            in1 => \N__13205\,
            in2 => \_gnd_net_\,
            in3 => \N__16795\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i9_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16792\,
            in1 => \N__14474\,
            in2 => \_gnd_net_\,
            in3 => \N__13273\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => \N__16686\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i1_3_lut_adj_117_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__16249\,
            in1 => \N__16778\,
            in2 => \_gnd_net_\,
            in3 => \N__13249\,
            lcout => n234,
            ltout => \n234_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.state_i1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011000000010"
        )
    port map (
            in0 => \N__15983\,
            in1 => \N__16187\,
            in2 => \N__13277\,
            in3 => \N__14089\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.writeByte_83_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__14090\,
            in1 => \N__15981\,
            in2 => \N__16198\,
            in3 => \N__16783\,
            lcout => \writeByte\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i10_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__16779\,
            in1 => \_gnd_net_\,
            in2 => \N__13274\,
            in3 => \N__16717\,
            lcout => \Inst_eia232.Inst_transmitter.txBuffer_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.state_i0_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__16031\,
            in1 => \N__15982\,
            in2 => \N__13259\,
            in3 => \N__16191\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i28_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__15980\,
            in1 => \N__14225\,
            in2 => \N__36422\,
            in3 => \N__21669\,
            lcout => \dataBuffer_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i25_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__21668\,
            in1 => \N__36402\,
            in2 => \N__13994\,
            in3 => \N__15984\,
            lcout => \dataBuffer_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byteDone_81_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001111"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__14108\,
            in2 => \N__16804\,
            in3 => \N__13343\,
            lcout => \byteDone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.bytes_i2_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__14180\,
            in1 => \N__14422\,
            in2 => \_gnd_net_\,
            in3 => \N__14146\,
            lcout => bytes_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37483\,
            ce => \N__13457\,
            sr => \N__13439\
        );

    \Inst_eia232.Inst_transmitter.bytes_i0_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__14147\,
            in1 => \_gnd_net_\,
            in2 => \N__14423\,
            in3 => \N__14178\,
            lcout => bytes_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37483\,
            ce => \N__13457\,
            sr => \N__13439\
        );

    \Inst_eia232.Inst_transmitter.bytes_i1_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14418\,
            lcout => bytes_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37483\,
            ce => \N__13457\,
            sr => \N__13439\
        );

    \Inst_eia232.Inst_transmitter.bits__i3_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__13379\,
            in1 => \N__13333\,
            in2 => \N__13370\,
            in3 => \N__13307\,
            lcout => \Inst_eia232.Inst_transmitter.bits_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => \N__13291\,
            sr => \N__16815\
        );

    \Inst_eia232.Inst_transmitter.bits__i2_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__13306\,
            in1 => \N__13365\,
            in2 => \_gnd_net_\,
            in3 => \N__13334\,
            lcout => \Inst_eia232.Inst_transmitter.bits_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => \N__13291\,
            sr => \N__16815\
        );

    \Inst_eia232.Inst_transmitter.i2_4_lut_adj_115_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__13412\,
            in1 => \N__13530\,
            in2 => \N__13480\,
            in3 => \N__13505\,
            lcout => n9,
            ltout => \n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i936_3_lut_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__16802\,
            in1 => \_gnd_net_\,
            in2 => \N__13382\,
            in3 => \N__13352\,
            lcout => n4082,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i2_4_lut_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__13378\,
            in1 => \N__13331\,
            in2 => \N__13369\,
            in3 => \N__13304\,
            lcout => n3493,
            ltout => \n3493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i5585_2_lut_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13346\,
            in3 => \N__16707\,
            lcout => n6749,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.bits__i1_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13332\,
            in2 => \_gnd_net_\,
            in3 => \N__13305\,
            lcout => \Inst_eia232.Inst_transmitter.bits_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => \N__13291\,
            sr => \N__16815\
        );

    \i1_2_lut_3_lut_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__16803\,
            in1 => \N__18505\,
            in2 => \_gnd_net_\,
            in3 => \N__16706\,
            lcout => n3615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.counter__i3_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__13410\,
            in1 => \N__13532\,
            in2 => \N__13481\,
            in3 => \N__13499\,
            lcout => \Inst_eia232.Inst_transmitter.counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37475\,
            ce => \N__13427\,
            sr => \N__16688\
        );

    \Inst_eia232.Inst_transmitter.i1166_2_lut_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13496\,
            in1 => \N__13407\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_transmitter.n2201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.counter__i4_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__13479\,
            in1 => \N__13531\,
            in2 => \N__13517\,
            in3 => \N__13514\,
            lcout => \Inst_eia232.Inst_transmitter.counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37475\,
            ce => \N__13427\,
            sr => \N__16688\
        );

    \Inst_eia232.Inst_transmitter.counter__i1_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__13497\,
            in1 => \N__13408\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_eia232.Inst_transmitter.counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37475\,
            ce => \N__13427\,
            sr => \N__16688\
        );

    \Inst_eia232.Inst_transmitter.i7274_2_lut_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13495\,
            in2 => \_gnd_net_\,
            in3 => \N__13513\,
            lcout => \Inst_eia232.Inst_transmitter.n8642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.counter__i2_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__13498\,
            in1 => \N__13409\,
            in2 => \_gnd_net_\,
            in3 => \N__13475\,
            lcout => \Inst_eia232.Inst_transmitter.counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37475\,
            ce => \N__13427\,
            sr => \N__16688\
        );

    \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_4_lut_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110010"
        )
    port map (
            in0 => \N__36346\,
            in1 => \N__15997\,
            in2 => \N__16070\,
            in3 => \N__16196\,
            lcout => \Inst_eia232.Inst_transmitter.n3594\,
            ltout => \Inst_eia232.Inst_transmitter.n3594_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i3560_2_lut_3_lut_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__16197\,
            in1 => \_gnd_net_\,
            in2 => \N__13442\,
            in3 => \N__15998\,
            lcout => \Inst_eia232.Inst_transmitter.n4719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.counter__i0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13411\,
            in2 => \_gnd_net_\,
            in3 => \N__13426\,
            lcout => \Inst_eia232.Inst_transmitter.counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37474\,
            ce => 'H',
            sr => \N__16687\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13601\,
            in2 => \_gnd_net_\,
            in3 => \N__36399\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37476\,
            ce => \N__21682\,
            sr => \N__15902\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i4_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__36401\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13589\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37476\,
            ce => \N__21682\,
            sr => \N__15902\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i5_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13580\,
            in2 => \_gnd_net_\,
            in3 => \N__36400\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37476\,
            ce => \N__21682\,
            sr => \N__15902\
        );

    \Inst_eia232.Inst_transmitter.txBuffer_i1_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13571\,
            lcout => tx_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37477\,
            ce => \N__16685\,
            sr => \N__16814\
        );

    \GENERIC_FIFO_1.write_pointer_919__i0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16616\,
            in2 => \_gnd_net_\,
            in3 => \N__13547\,
            lcout => \GENERIC_FIFO_1.write_pointer_0\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \GENERIC_FIFO_1.n7836\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16568\,
            in2 => \_gnd_net_\,
            in3 => \N__13544\,
            lcout => \GENERIC_FIFO_1.write_pointer_1\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7836\,
            carryout => \GENERIC_FIFO_1.n7837\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16516\,
            in2 => \_gnd_net_\,
            in3 => \N__13541\,
            lcout => \GENERIC_FIFO_1.write_pointer_2\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7837\,
            carryout => \GENERIC_FIFO_1.n7838\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i3_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16469\,
            in2 => \_gnd_net_\,
            in3 => \N__13538\,
            lcout => \GENERIC_FIFO_1.write_pointer_3\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7838\,
            carryout => \GENERIC_FIFO_1.n7839\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i4_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14934\,
            in2 => \_gnd_net_\,
            in3 => \N__13535\,
            lcout => \GENERIC_FIFO_1.write_pointer_4\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7839\,
            carryout => \GENERIC_FIFO_1.n7840\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i5_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14863\,
            in2 => \_gnd_net_\,
            in3 => \N__13625\,
            lcout => \GENERIC_FIFO_1.write_pointer_5\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7840\,
            carryout => \GENERIC_FIFO_1.n7841\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i6_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17102\,
            in2 => \_gnd_net_\,
            in3 => \N__13622\,
            lcout => \GENERIC_FIFO_1.write_pointer_6\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7841\,
            carryout => \GENERIC_FIFO_1.n7842\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i7_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14567\,
            in2 => \_gnd_net_\,
            in3 => \N__13619\,
            lcout => \GENERIC_FIFO_1.write_pointer_7\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7842\,
            carryout => \GENERIC_FIFO_1.n7843\,
            clk => \N__37482\,
            ce => \N__14981\,
            sr => \N__14822\
        );

    \GENERIC_FIFO_1.write_pointer_919__i8_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14657\,
            in2 => \_gnd_net_\,
            in3 => \N__13616\,
            lcout => \GENERIC_FIFO_1.write_pointer_8\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \GENERIC_FIFO_1.n7844\,
            clk => \N__37489\,
            ce => \N__14996\,
            sr => \N__14821\
        );

    \GENERIC_FIFO_1.write_pointer_919__i9_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14611\,
            in2 => \_gnd_net_\,
            in3 => \N__13613\,
            lcout => \GENERIC_FIFO_1.write_pointer_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37489\,
            ce => \N__14996\,
            sr => \N__14821\
        );

    \GENERIC_FIFO_1.add_6561_2_lut_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14792\,
            in2 => \N__13814\,
            in3 => \_gnd_net_\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_0\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \GENERIC_FIFO_1.n7827\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_3_lut_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13802\,
            in2 => \N__14786\,
            in3 => \N__13610\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_1\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7827\,
            carryout => \GENERIC_FIFO_1.n7828\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_4_lut_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13790\,
            in2 => \N__15092\,
            in3 => \N__13607\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_2\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7828\,
            carryout => \GENERIC_FIFO_1.n7829\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_5_lut_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13778\,
            in2 => \N__15080\,
            in3 => \N__13604\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_3\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7829\,
            carryout => \GENERIC_FIFO_1.n7830\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_6_lut_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13766\,
            in2 => \N__15068\,
            in3 => \N__13700\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_4\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7830\,
            carryout => \GENERIC_FIFO_1.n7831\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_7_lut_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13751\,
            in2 => \N__15056\,
            in3 => \N__13697\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_5\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7831\,
            carryout => \GENERIC_FIFO_1.n7832\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_8_lut_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13739\,
            in2 => \N__15044\,
            in3 => \N__13694\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_6\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7832\,
            carryout => \GENERIC_FIFO_1.n7833\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_9_lut_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13727\,
            in2 => \N__15029\,
            in3 => \N__13691\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_7\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7833\,
            carryout => \GENERIC_FIFO_1.n7834\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_10_lut_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15017\,
            in2 => \N__13715\,
            in3 => \N__13688\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_8\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \GENERIC_FIFO_1.n7835\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_6561_11_lut_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13826\,
            in1 => \N__15005\,
            in2 => \_gnd_net_\,
            in3 => \N__13685\,
            lcout => \GENERIC_FIFO_1.level_9_N_876_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i7_4_lut_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13681\,
            in1 => \N__13667\,
            in2 => \N__13655\,
            in3 => \N__13637\,
            lcout => \GENERIC_FIFO_1.n17_adj_1278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i6_1_lut_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14868\,
            lcout => \GENERIC_FIFO_1.n1375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i7282_4_lut_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13682\,
            in1 => \N__13666\,
            in2 => \N__13654\,
            in3 => \N__13636\,
            lcout => \GENERIC_FIFO_1.n8650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_2_lut_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17233\,
            in2 => \N__16630\,
            in3 => \_gnd_net_\,
            lcout => \GENERIC_FIFO_1.n12\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \GENERIC_FIFO_1.n7818\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_3_lut_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16575\,
            in2 => \_gnd_net_\,
            in3 => \N__13793\,
            lcout => \GENERIC_FIFO_1.n11\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7818\,
            carryout => \GENERIC_FIFO_1.n7819\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_4_lut_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16531\,
            in2 => \_gnd_net_\,
            in3 => \N__13781\,
            lcout => \GENERIC_FIFO_1.n10\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7819\,
            carryout => \GENERIC_FIFO_1.n7820\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_5_lut_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16483\,
            in2 => \_gnd_net_\,
            in3 => \N__13769\,
            lcout => \GENERIC_FIFO_1.n9\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7820\,
            carryout => \GENERIC_FIFO_1.n7821\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_6_lut_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14938\,
            in2 => \_gnd_net_\,
            in3 => \N__13754\,
            lcout => \GENERIC_FIFO_1.n8\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7821\,
            carryout => \GENERIC_FIFO_1.n7822\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_7_lut_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14875\,
            in2 => \_gnd_net_\,
            in3 => \N__13742\,
            lcout => \GENERIC_FIFO_1.n7\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7822\,
            carryout => \GENERIC_FIFO_1.n7823\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_8_lut_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17116\,
            in2 => \_gnd_net_\,
            in3 => \N__13730\,
            lcout => \GENERIC_FIFO_1.n6\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7823\,
            carryout => \GENERIC_FIFO_1.n7824\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_9_lut_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14572\,
            in2 => \_gnd_net_\,
            in3 => \N__13718\,
            lcout => \GENERIC_FIFO_1.n5\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7824\,
            carryout => \GENERIC_FIFO_1.n7825\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_10_lut_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14662\,
            in2 => \_gnd_net_\,
            in3 => \N__13703\,
            lcout => \GENERIC_FIFO_1.n4\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \GENERIC_FIFO_1.n7826\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_1_11_lut_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14616\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13829\,
            lcout => \GENERIC_FIFO_1.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i9_1_lut_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14661\,
            lcout => \GENERIC_FIFO_1.n1372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i8_1_lut_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14571\,
            lcout => \GENERIC_FIFO_1.n1373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i10_1_lut_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14615\,
            lcout => \GENERIC_FIFO_1.n1371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i8_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36413\,
            in2 => \_gnd_net_\,
            in3 => \N__15999\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37527\,
            ce => \N__21655\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i20_3_lut_3_lut_4_lut_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110010"
        )
    port map (
            in0 => \N__36406\,
            in1 => \N__15985\,
            in2 => \N__16069\,
            in3 => \N__16192\,
            lcout => n4005,
            ltout => \n4005_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i14_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__15986\,
            in1 => \N__13841\,
            in2 => \N__13817\,
            in3 => \N__36410\,
            lcout => \dataBuffer_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i22_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__36408\,
            in1 => \N__13931\,
            in2 => \N__21657\,
            in3 => \N__15991\,
            lcout => \dataBuffer_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i24_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__15988\,
            in1 => \N__21611\,
            in2 => \N__13913\,
            in3 => \N__36412\,
            lcout => \dataBuffer_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i19_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__36407\,
            in1 => \N__13861\,
            in2 => \N__21656\,
            in3 => \N__15990\,
            lcout => \dataBuffer_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i18_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__15987\,
            in1 => \N__21610\,
            in2 => \N__14033\,
            in3 => \N__36411\,
            lcout => \dataBuffer_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.mux_650_i7_3_lut_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13921\,
            in1 => \N__13930\,
            in2 => \_gnd_net_\,
            in3 => \N__13960\,
            lcout => \Inst_eia232.Inst_transmitter.n1323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i30_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__15989\,
            in1 => \N__36409\,
            in2 => \N__21658\,
            in3 => \N__13922\,
            lcout => \dataBuffer_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byte__i0_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__14749\,
            in1 => \N__13912\,
            in2 => \N__13964\,
            in3 => \N__13868\,
            lcout => \Inst_eia232.Inst_transmitter.byte_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => \N__14075\,
            sr => \N__16232\
        );

    \Inst_eia232.Inst_transmitter.i2444_3_lut_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13889\,
            in1 => \N__13880\,
            in2 => \_gnd_net_\,
            in3 => \N__16128\,
            lcout => \Inst_eia232.Inst_transmitter.n3571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i7532_2_lut_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16130\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14303\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_transmitter.n8854_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byte__i3_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__13959\,
            in1 => \N__13862\,
            in2 => \N__13850\,
            in3 => \N__14751\,
            lcout => \Inst_eia232.Inst_transmitter.byte_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => \N__14075\,
            sr => \N__16232\
        );

    \Inst_eia232.Inst_transmitter.i2505_3_lut_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16131\,
            in1 => \N__13840\,
            in2 => \_gnd_net_\,
            in3 => \N__14276\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_transmitter.n3632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byte__i6_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14048\,
            in2 => \N__14042\,
            in3 => \N__14752\,
            lcout => \Inst_eia232.Inst_transmitter.byte_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => \N__14075\,
            sr => \N__16232\
        );

    \Inst_eia232.Inst_transmitter.i7530_2_lut_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16129\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14333\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_transmitter.n8851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byte__i2_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__13958\,
            in1 => \N__14032\,
            in2 => \N__14018\,
            in3 => \N__14750\,
            lcout => \Inst_eia232.Inst_transmitter.byte_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => \N__14075\,
            sr => \N__16232\
        );

    \Inst_eia232.Inst_transmitter.byte__i1_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__13979\,
            in1 => \N__14753\,
            in2 => \N__16132\,
            in3 => \N__14362\,
            lcout => \Inst_eia232.Inst_transmitter.byte_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37498\,
            ce => \N__14071\,
            sr => \N__16228\
        );

    \Inst_eia232.Inst_transmitter.i3105_2_lut_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15951\,
            in2 => \_gnd_net_\,
            in3 => \N__16173\,
            lcout => n4248,
            ltout => \n4248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_130_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__14416\,
            in1 => \N__14144\,
            in2 => \N__14000\,
            in3 => \N__14176\,
            lcout => n1336,
            ltout => \n1336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i5539_2_lut_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13997\,
            in3 => \N__14059\,
            lcout => \Inst_eia232.Inst_transmitter.n6703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i7569_2_lut_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13990\,
            in2 => \_gnd_net_\,
            in3 => \N__13957\,
            lcout => \Inst_eia232.Inst_transmitter.n8847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010000000"
        )
    port map (
            in0 => \N__14177\,
            in1 => \N__14417\,
            in2 => \N__13973\,
            in3 => \N__14145\,
            lcout => n1320,
            ltout => \n1320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i7548_2_lut_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14228\,
            in3 => \N__14224\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_transmitter.n8756_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byte__i4_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__14754\,
            in1 => \N__16121\,
            in2 => \N__14213\,
            in3 => \N__14210\,
            lcout => \Inst_eia232.Inst_transmitter.byte_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37498\,
            ce => \N__14071\,
            sr => \N__16228\
        );

    \i7565_3_lut_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__14142\,
            in1 => \N__14412\,
            in2 => \_gnd_net_\,
            in3 => \N__14173\,
            lcout => \state_1_N_371_1\,
            ltout => \state_1_N_371_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i5581_2_lut_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__16178\,
            in1 => \_gnd_net_\,
            in2 => \N__14189\,
            in3 => \_gnd_net_\,
            lcout => \Inst_eia232.Inst_transmitter.n6745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.bytes_2__I_0_i3_3_lut_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14501\,
            in1 => \N__14186\,
            in2 => \_gnd_net_\,
            in3 => \N__14174\,
            lcout => \Inst_eia232.Inst_transmitter.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.bytes_2__I_0_i1_3_lut_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14413\,
            in1 => \N__14260\,
            in2 => \_gnd_net_\,
            in3 => \N__21539\,
            lcout => \Inst_eia232.Inst_transmitter.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i1201_rep_51_2_lut_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14415\,
            in2 => \_gnd_net_\,
            in3 => \N__14175\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_transmitter.n9218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.disabled_90_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__14239\,
            in1 => \N__14143\,
            in2 => \N__14117\,
            in3 => \N__14114\,
            lcout => disabled,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37492\,
            ce => \N__14099\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i1_3_lut_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__15967\,
            in1 => \N__16177\,
            in2 => \_gnd_net_\,
            in3 => \N__14088\,
            lcout => \Inst_eia232.Inst_transmitter.n3652\,
            ltout => \Inst_eia232.Inst_transmitter.n3652_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i2_3_lut_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__14414\,
            in1 => \_gnd_net_\,
            in2 => \N__14384\,
            in3 => \N__14381\,
            lcout => \Inst_eia232.Inst_transmitter.n2580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i1_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__14375\,
            in1 => \N__21732\,
            in2 => \N__14363\,
            in3 => \N__21664\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i2_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__21662\,
            in1 => \N__14345\,
            in2 => \N__21742\,
            in3 => \N__14332\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i3_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__14302\,
            in1 => \N__21733\,
            in2 => \N__14318\,
            in3 => \N__21665\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i6_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__21663\,
            in1 => \N__14288\,
            in2 => \N__21743\,
            in3 => \N__14275\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.disabledBuffer_i1_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__14249\,
            in1 => \N__21741\,
            in2 => \N__21676\,
            in3 => \N__14261\,
            lcout => \Inst_eia232.Inst_transmitter.disabledBuffer_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.disabledGroupsReg_i0_i1_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22291\,
            in1 => \N__26730\,
            in2 => \_gnd_net_\,
            in3 => \N__14248\,
            lcout => \disabledGroupsReg_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.disabledBuffer_i3_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__14240\,
            in1 => \N__21734\,
            in2 => \N__21677\,
            in3 => \N__14510\,
            lcout => \Inst_eia232.Inst_transmitter.disabledBuffer_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.disabledGroupsReg_i0_i3_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14509\,
            in1 => \_gnd_net_\,
            in2 => \N__22295\,
            in3 => \N__31398\,
            lcout => \disabledGroupsReg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.disabledBuffer_i2_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__21729\,
            in1 => \N__14500\,
            in2 => \N__14486\,
            in3 => \N__21667\,
            lcout => \Inst_eia232.Inst_transmitter.disabledBuffer_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.disabledGroupsReg_i0_i2_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22277\,
            in1 => \N__29127\,
            in2 => \_gnd_net_\,
            in3 => \N__14482\,
            lcout => \disabledGroupsReg_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byte__i7_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__14467\,
            in1 => \N__14758\,
            in2 => \N__14444\,
            in3 => \N__16091\,
            lcout => \Inst_eia232.Inst_transmitter.byte_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i5_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21889\,
            in1 => \N__31406\,
            in2 => \_gnd_net_\,
            in3 => \N__14773\,
            lcout => \maskRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register_80_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100010001"
        )
    port map (
            in0 => \N__15695\,
            in1 => \N__14888\,
            in2 => \_gnd_net_\,
            in3 => \N__26291\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_6_i1_1_lut_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17057\,
            lcout => \GENERIC_FIFO_1.level_9_N_925_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.dataBuffer_i7_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21666\,
            in1 => \N__14456\,
            in2 => \N__14443\,
            in3 => \N__21730\,
            lcout => \Inst_eia232.Inst_transmitter.dataBuffer_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_2_lut_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16346\,
            in1 => \N__17065\,
            in2 => \_gnd_net_\,
            in3 => \N__14429\,
            lcout => \GENERIC_FIFO_1.n8779\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \GENERIC_FIFO_1.n7929\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_3_lut_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16343\,
            in1 => \N__19415\,
            in2 => \_gnd_net_\,
            in3 => \N__14426\,
            lcout => \GENERIC_FIFO_1.n8813\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7929\,
            carryout => \GENERIC_FIFO_1.n7930\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_4_lut_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16349\,
            in1 => \N__19343\,
            in2 => \_gnd_net_\,
            in3 => \N__14534\,
            lcout => \GENERIC_FIFO_1.n8814\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7930\,
            carryout => \GENERIC_FIFO_1.n7931\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_5_lut_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16341\,
            in1 => \N__18980\,
            in2 => \_gnd_net_\,
            in3 => \N__14531\,
            lcout => \GENERIC_FIFO_1.n8815\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7931\,
            carryout => \GENERIC_FIFO_1.n7932\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_6_lut_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16347\,
            in1 => \N__19259\,
            in2 => \_gnd_net_\,
            in3 => \N__14528\,
            lcout => \GENERIC_FIFO_1.n8816\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7932\,
            carryout => \GENERIC_FIFO_1.n7933\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_7_lut_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16342\,
            in1 => \N__19190\,
            in2 => \_gnd_net_\,
            in3 => \N__14525\,
            lcout => \GENERIC_FIFO_1.n8817\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7933\,
            carryout => \GENERIC_FIFO_1.n7934\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_8_lut_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16348\,
            in1 => \N__19118\,
            in2 => \_gnd_net_\,
            in3 => \N__14522\,
            lcout => \GENERIC_FIFO_1.n8818\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7934\,
            carryout => \GENERIC_FIFO_1.n7935\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_9_lut_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16340\,
            in1 => \N__19757\,
            in2 => \_gnd_net_\,
            in3 => \N__14519\,
            lcout => \GENERIC_FIFO_1.n8819\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7935\,
            carryout => \GENERIC_FIFO_1.n7936\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_10_lut_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16345\,
            in1 => \N__19565\,
            in2 => \_gnd_net_\,
            in3 => \N__14516\,
            lcout => \GENERIC_FIFO_1.n8820\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \GENERIC_FIFO_1.n7937\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_add_4_11_lut_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16344\,
            in1 => \N__17177\,
            in2 => \_gnd_net_\,
            in3 => \N__14513\,
            lcout => \GENERIC_FIFO_1.n8821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105_bdd_4_lut_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__25500\,
            in1 => \N__22074\,
            in2 => \N__28086\,
            in3 => \N__14810\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3584_1_lut_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14774\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.byte__i5_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__14701\,
            in1 => \N__14759\,
            in2 => \N__14717\,
            in3 => \N__16087\,
            lcout => \Inst_eia232.Inst_transmitter.byte_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i7308_3_lut_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__16976\,
            in1 => \N__16925\,
            in2 => \_gnd_net_\,
            in3 => \N__17255\,
            lcout => OPEN,
            ltout => \GENERIC_FIFO_1.n8677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i1_4_lut_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__17306\,
            in1 => \N__16877\,
            in2 => \N__14690\,
            in3 => \N__17234\,
            lcout => \GENERIC_FIFO_1.n1396\,
            ltout => \GENERIC_FIFO_1.n1396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i2_4_lut_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__36644\,
            in1 => \N__30154\,
            in2 => \N__14687\,
            in3 => \N__15269\,
            lcout => \GENERIC_FIFO_1.fifo_memory_N_983\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i5_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__15827\,
            in1 => \N__20580\,
            in2 => \N__18695\,
            in3 => \N__25512\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37484\,
            ce => 'H',
            sr => \N__14684\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110010101101010"
        )
    port map (
            in0 => \N__20309\,
            in1 => \N__20798\,
            in2 => \N__30357\,
            in3 => \N__31816\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37491\,
            ce => 'H',
            sr => \N__18791\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22415\,
            in1 => \N__29789\,
            in2 => \N__26831\,
            in3 => \N__14678\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i7_4_lut_adj_122_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14930\,
            in1 => \N__14656\,
            in2 => \N__14617\,
            in3 => \N__14566\,
            lcout => OPEN,
            ltout => \GENERIC_FIFO_1.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i9_4_lut_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17101\,
            in1 => \N__16468\,
            in2 => \N__14999\,
            in3 => \N__14971\,
            lcout => \GENERIC_FIFO_1.n20_adj_1274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i5_1_lut_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14929\,
            lcout => \GENERIC_FIFO_1.n1376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i4_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111011010010"
        )
    port map (
            in0 => \N__28087\,
            in1 => \N__20598\,
            in2 => \N__19070\,
            in3 => \N__15851\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37497\,
            ce => 'H',
            sr => \N__18860\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_adj_70_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14903\,
            in1 => \N__14897\,
            in2 => \N__16862\,
            in3 => \N__15212\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i5_2_lut_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16567\,
            in2 => \_gnd_net_\,
            in3 => \N__16615\,
            lcout => OPEN,
            ltout => \GENERIC_FIFO_1.n16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i10_4_lut_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14864\,
            in1 => \N__16517\,
            in2 => \N__14831\,
            in3 => \N__14828\,
            lcout => \GENERIC_FIFO_1.n4721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_7715_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__23038\,
            in1 => \N__30432\,
            in2 => \N__22087\,
            in3 => \N__22172\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_2_lut_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14801\,
            in2 => \N__15239\,
            in3 => \_gnd_net_\,
            lcout => \GENERIC_FIFO_1.n24\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \GENERIC_FIFO_1.n7809\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_3_lut_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19466\,
            in2 => \_gnd_net_\,
            in3 => \N__14777\,
            lcout => \GENERIC_FIFO_1.n23\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7809\,
            carryout => \GENERIC_FIFO_1.n7810\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_4_lut_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16832\,
            in2 => \_gnd_net_\,
            in3 => \N__15083\,
            lcout => \GENERIC_FIFO_1.n22\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7810\,
            carryout => \GENERIC_FIFO_1.n7811\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_5_lut_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19049\,
            in2 => \_gnd_net_\,
            in3 => \N__15071\,
            lcout => \GENERIC_FIFO_1.n21\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7811\,
            carryout => \GENERIC_FIFO_1.n7812\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_6_lut_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16841\,
            in2 => \_gnd_net_\,
            in3 => \N__15059\,
            lcout => \GENERIC_FIFO_1.n20\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7812\,
            carryout => \GENERIC_FIFO_1.n7813\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_7_lut_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16379\,
            in2 => \_gnd_net_\,
            in3 => \N__15047\,
            lcout => \GENERIC_FIFO_1.n19\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7813\,
            carryout => \GENERIC_FIFO_1.n7814\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_8_lut_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19454\,
            in2 => \_gnd_net_\,
            in3 => \N__15032\,
            lcout => \GENERIC_FIFO_1.n18_adj_1275\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7814\,
            carryout => \GENERIC_FIFO_1.n7815\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_9_lut_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15218\,
            in2 => \_gnd_net_\,
            in3 => \N__15020\,
            lcout => \GENERIC_FIFO_1.n17\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7815\,
            carryout => \GENERIC_FIFO_1.n7816\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_10_lut_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19298\,
            in2 => \_gnd_net_\,
            in3 => \N__15011\,
            lcout => \GENERIC_FIFO_1.n16_adj_1273\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \GENERIC_FIFO_1.n7817\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_912_1372_add_1_add_2_11_lut_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17132\,
            in2 => \_gnd_net_\,
            in3 => \N__15008\,
            lcout => \GENERIC_FIFO_1.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i7312_4_lut_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15136\,
            in1 => \N__15121\,
            in2 => \N__15230\,
            in3 => \N__15275\,
            lcout => \GENERIC_FIFO_1.n8681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i1_3_lut_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15736\,
            in1 => \N__17069\,
            in2 => \_gnd_net_\,
            in3 => \N__19612\,
            lcout => \GENERIC_FIFO_1.n78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i680_1_lut_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17229\,
            lcout => \GENERIC_FIFO_1.level_9__N_900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i7286_4_lut_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15151\,
            in1 => \N__15163\,
            in2 => \N__15188\,
            in3 => \N__15199\,
            lcout => \GENERIC_FIFO_1.n8654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i8_1_lut_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19752\,
            lcout => \GENERIC_FIFO_1.n1418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i6_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101100101101010"
        )
    port map (
            in0 => \N__18758\,
            in1 => \N__20603\,
            in2 => \N__15803\,
            in3 => \N__30461\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37526\,
            ce => 'H',
            sr => \N__18836\
        );

    \GENERIC_FIFO_1.i6_4_lut_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15203\,
            in1 => \N__15187\,
            in2 => \N__15170\,
            in3 => \N__15152\,
            lcout => OPEN,
            ltout => \GENERIC_FIFO_1.n16_adj_1276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i8_3_lut_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15140\,
            in2 => \N__15125\,
            in3 => \N__15122\,
            lcout => \GENERIC_FIFO_1.n18_adj_1277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i1_4_lut_adj_119_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__15110\,
            in1 => \N__36414\,
            in2 => \N__15104\,
            in3 => \N__15371\,
            lcout => \GENERIC_FIFO_1.n141\,
            ltout => \GENERIC_FIFO_1.n141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i10_3_lut_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17176\,
            in2 => \N__15365\,
            in3 => \N__17194\,
            lcout => \GENERIC_FIFO_1.n69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_prescaler.counter_922_923__i2_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18553\,
            lcout => \Inst_eia232.Inst_prescaler.counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37538\,
            ce => 'H',
            sr => \N__18434\
        );

    \Inst_eia232.Inst_prescaler.counter_922_923__i1_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18527\,
            lcout => \Inst_eia232.Inst_prescaler.counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37538\,
            ce => 'H',
            sr => \N__18434\
        );

    \Inst_eia232.Inst_receiver.bitcount_i2_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001011110000"
        )
    port map (
            in0 => \N__15293\,
            in1 => \N__20185\,
            in2 => \N__15320\,
            in3 => \N__15337\,
            lcout => \Inst_eia232.Inst_receiver.bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \N__17717\
        );

    \Inst_eia232.Inst_receiver.i1108_2_lut_3_lut_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__20182\,
            in1 => \_gnd_net_\,
            in2 => \N__15338\,
            in3 => \N__15290\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n2143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.bitcount_i3_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__15319\,
            in1 => \_gnd_net_\,
            in2 => \N__15341\,
            in3 => \N__15304\,
            lcout => \Inst_eia232.Inst_receiver.bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \N__17717\
        );

    \Inst_eia232.Inst_receiver.bitcount_i0_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__20183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15291\,
            lcout => \Inst_eia232.Inst_receiver.bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \N__17717\
        );

    \Inst_eia232.Inst_receiver.bitcount_i1_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__15292\,
            in1 => \N__20184\,
            in2 => \_gnd_net_\,
            in3 => \N__15336\,
            lcout => \Inst_eia232.Inst_receiver.bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \N__17717\
        );

    \Inst_eia232.Inst_receiver.i3_4_lut_adj_79_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__15332\,
            in1 => \N__15315\,
            in2 => \N__15305\,
            in3 => \N__15289\,
            lcout => \Inst_eia232.Inst_receiver.n7_adj_1264\,
            ltout => \Inst_eia232.Inst_receiver.n7_adj_1264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7493_4_lut_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__15397\,
            in1 => \N__20181\,
            in2 => \N__15428\,
            in3 => \N__15419\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n8769_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i24_4_lut_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000110001"
        )
    port map (
            in0 => \N__17861\,
            in1 => \N__17935\,
            in2 => \N__15425\,
            in3 => \N__17674\,
            lcout => n3753,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_4_lut_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__20134\,
            in1 => \N__15511\,
            in2 => \N__15398\,
            in3 => \N__15412\,
            lcout => \Inst_eia232.Inst_receiver.n5504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.bytecount_i1_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010011100"
        )
    port map (
            in0 => \N__20164\,
            in1 => \N__15395\,
            in2 => \N__20135\,
            in3 => \N__20211\,
            lcout => \Inst_eia232.Inst_receiver.bytecount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37540\,
            ce => \N__20098\,
            sr => \N__16274\
        );

    \Inst_eia232.Inst_receiver.i5572_2_lut_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20129\,
            in2 => \_gnd_net_\,
            in3 => \N__20163\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n6736_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.bytecount_i2_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__15413\,
            in1 => \N__15396\,
            in2 => \N__15422\,
            in3 => \N__20212\,
            lcout => \Inst_eia232.Inst_receiver.bytecount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37540\,
            ce => \N__20098\,
            sr => \N__16274\
        );

    \Inst_eia232.Inst_receiver.i7495_2_lut_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20128\,
            in2 => \_gnd_net_\,
            in3 => \N__15410\,
            lcout => \Inst_eia232.Inst_receiver.n8772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7214_2_lut_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15411\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15391\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n8582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7549_4_lut_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__20133\,
            in1 => \N__20209\,
            in2 => \N__15374\,
            in3 => \N__20162\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n8831_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i25_4_lut_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001010001"
        )
    port map (
            in0 => \N__17976\,
            in1 => \N__17862\,
            in2 => \N__15443\,
            in3 => \N__17673\,
            lcout => \Inst_eia232.Inst_receiver.n3718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i7_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15509\,
            in1 => \N__34774\,
            in2 => \N__15550\,
            in3 => \N__18228\,
            lcout => cmd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i6_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__18226\,
            in1 => \N__15545\,
            in2 => \N__18375\,
            in3 => \N__34809\,
            lcout => \Inst_eia232.Inst_receiver.cmd_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_98_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__15508\,
            in1 => \N__18364\,
            in2 => \N__15549\,
            in3 => \N__18408\,
            lcout => \Inst_eia232.Inst_receiver.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_97_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__18363\,
            in1 => \N__15538\,
            in2 => \N__18415\,
            in3 => \N__15506\,
            lcout => \Inst_eia232.Inst_receiver.n14_adj_1265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i8_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__15510\,
            in1 => \N__34773\,
            in2 => \N__18484\,
            in3 => \N__18229\,
            lcout => \nstate_2_N_241_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15537\,
            in2 => \_gnd_net_\,
            in3 => \N__15507\,
            lcout => \Inst_eia232.Inst_receiver.n5498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i4_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__18414\,
            in1 => \N__18060\,
            in2 => \N__34839\,
            in3 => \N__18227\,
            lcout => \Inst_eia232.Inst_receiver.cmd_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i5_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__18225\,
            in1 => \N__34805\,
            in2 => \N__18376\,
            in3 => \N__18413\,
            lcout => \Inst_eia232.Inst_receiver.cmd_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i1_2_lut_adj_114_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15475\,
            in2 => \_gnd_net_\,
            in3 => \N__15452\,
            lcout => \Inst_eia232.Inst_transmitter.n3552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.xon_33_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__18310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15461\,
            lcout => \Inst_eia232.xon\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37518\,
            ce => 'H',
            sr => \N__17487\
        );

    \Inst_core.Inst_decoder.wrtrigcfg__i2_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18058\,
            in1 => \N__18131\,
            in2 => \N__18203\,
            in3 => \N__15586\,
            lcout => wrtrigcfg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37518\,
            ce => 'H',
            sr => \N__17487\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_94_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__18129\,
            in1 => \N__18193\,
            in2 => \_gnd_net_\,
            in3 => \N__18057\,
            lcout => \Inst_eia232.Inst_receiver.n75\,
            ltout => \Inst_eia232.Inst_receiver.n75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i2_4_lut_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__18412\,
            in1 => \N__18374\,
            in2 => \N__15464\,
            in3 => \N__15562\,
            lcout => \Inst_eia232.Inst_receiver.n5597\,
            ltout => \Inst_eia232.Inst_receiver.n5597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.xoff_34_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__18309\,
            in1 => \_gnd_net_\,
            in2 => \N__15455\,
            in3 => \_gnd_net_\,
            lcout => \Inst_eia232.xoff\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37518\,
            ce => 'H',
            sr => \N__17487\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_adj_84_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18308\,
            in2 => \_gnd_net_\,
            in3 => \N__15631\,
            lcout => \Inst_eia232.Inst_receiver.n90\,
            ltout => \Inst_eia232.Inst_receiver.n90_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_decoder.wrtrigcfg__i1_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18130\,
            in1 => \N__18194\,
            in2 => \N__15446\,
            in3 => \N__18059\,
            lcout => wrtrigcfg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37518\,
            ce => 'H',
            sr => \N__17487\
        );

    \Inst_core.Inst_decoder.wrtrigval__i0_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__15634\,
            in1 => \N__18295\,
            in2 => \_gnd_net_\,
            in3 => \N__17522\,
            lcout => wrtrigval_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => 'H',
            sr => \N__17494\
        );

    \Inst_eia232.id_32_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__18008\,
            in1 => \N__18339\,
            in2 => \N__18316\,
            in3 => \N__15572\,
            lcout => \Inst_eia232.id\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => 'H',
            sr => \N__17494\
        );

    \Inst_core.Inst_decoder.reset_52_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15571\,
            in1 => \N__18340\,
            in2 => \N__18017\,
            in3 => \N__18302\,
            lcout => \Inst_core.resetCmd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => 'H',
            sr => \N__17494\
        );

    \Inst_core.Inst_decoder.arm_53_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__17521\,
            in1 => \N__18338\,
            in2 => \N__18317\,
            in3 => \N__15570\,
            lcout => \Inst_core.arm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => 'H',
            sr => \N__17494\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_adj_81_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18293\,
            in2 => \_gnd_net_\,
            in3 => \N__18006\,
            lcout => OPEN,
            ltout => \n5698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_decoder.wrFlags_35_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18341\,
            in1 => \N__15551\,
            in2 => \N__15518\,
            in3 => \N__15515\,
            lcout => \wrFlags\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => 'H',
            sr => \N__17494\
        );

    \Inst_core.Inst_decoder.wrtrigmask__i0_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15635\,
            in1 => \N__18294\,
            in2 => \_gnd_net_\,
            in3 => \N__18009\,
            lcout => wrtrigmask_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => 'H',
            sr => \N__17494\
        );

    \Inst_core.Inst_decoder.wrtrigcfg__i0_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__18007\,
            in1 => \N__18307\,
            in2 => \_gnd_net_\,
            in3 => \N__15633\,
            lcout => wrtrigcfg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => 'H',
            sr => \N__17494\
        );

    \Inst_core.Inst_decoder.wrtrigval__i2_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__15608\,
            in1 => \N__18073\,
            in2 => \N__18200\,
            in3 => \N__18127\,
            lcout => wrtrigval_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \N__17495\
        );

    \Inst_core.Inst_decoder.wrtrigmask__i3_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18126\,
            in1 => \N__18179\,
            in2 => \N__18082\,
            in3 => \N__15604\,
            lcout => wrtrigmask_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \N__17495\
        );

    \Inst_core.Inst_decoder.wrtrigval__i1_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15605\,
            in1 => \N__18074\,
            in2 => \N__18201\,
            in3 => \N__18122\,
            lcout => wrtrigval_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \N__17495\
        );

    \Inst_core.Inst_decoder.wrtrigmask__i1_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__18124\,
            in1 => \N__18178\,
            in2 => \N__18081\,
            in3 => \N__15606\,
            lcout => wrtrigmask_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \N__17495\
        );

    \Inst_core.Inst_decoder.wrtrigmask__i2_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__15607\,
            in1 => \N__18069\,
            in2 => \N__18199\,
            in3 => \N__18125\,
            lcout => wrtrigmask_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \N__17495\
        );

    \Inst_eia232.Inst_receiver.i132_2_lut_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18289\,
            in2 => \_gnd_net_\,
            in3 => \N__15632\,
            lcout => \Inst_eia232.Inst_receiver.n112\,
            ltout => \Inst_eia232.Inst_receiver.n112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_decoder.wrtrigval__i3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__18177\,
            in1 => \N__18075\,
            in2 => \N__15590\,
            in3 => \N__18128\,
            lcout => wrtrigval_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \N__17495\
        );

    \Inst_core.Inst_decoder.wrtrigcfg__i3_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18123\,
            in1 => \N__15587\,
            in2 => \N__18083\,
            in3 => \N__18189\,
            lcout => wrtrigcfg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \N__17495\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i7_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__34356\,
            in1 => \N__34820\,
            in2 => \N__27208\,
            in3 => \N__34935\,
            lcout => cmd_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i7_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27023\,
            in1 => \N__27193\,
            in2 => \_gnd_net_\,
            in3 => \N__26470\,
            lcout => \maskRegister_7_adj_1321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i0_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35956\,
            in1 => \_gnd_net_\,
            in2 => \N__20690\,
            in3 => \N__15718\,
            lcout => \valueRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i31_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24049\,
            in1 => \N__34819\,
            in2 => \N__20447\,
            in3 => \N__34934\,
            lcout => cmd_38,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_flags.demux_15_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35955\,
            in1 => \N__22256\,
            in2 => \_gnd_net_\,
            in3 => \N__26244\,
            lcout => \flagDemux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i0_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15740\,
            in1 => \N__17052\,
            in2 => \_gnd_net_\,
            in3 => \N__19706\,
            lcout => \GENERIC_FIFO_1.read_pointer_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__15872\,
            in1 => \N__15719\,
            in2 => \N__20602\,
            in3 => \N__31796\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37481\,
            ce => 'H',
            sr => \N__20423\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__30936\,
            in1 => \N__32353\,
            in2 => \N__22088\,
            in3 => \N__22171\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_bdd_4_lut_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__33653\,
            in1 => \N__31795\,
            in2 => \N__15707\,
            in3 => \N__22086\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n9114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_762_i1_3_lut_4_lut_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__21911\,
            in1 => \N__15668\,
            in2 => \N__15704\,
            in3 => \N__24118\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18584\,
            in1 => \N__20519\,
            in2 => \N__18614\,
            in3 => \N__15701\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_706_i1_3_lut_4_lut_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__21910\,
            in1 => \N__15655\,
            in2 => \N__15683\,
            in3 => \N__24119\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__26270\,
            in1 => \N__15667\,
            in2 => \N__15656\,
            in3 => \N__18677\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i1_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15651\,
            in1 => \N__15864\,
            in2 => \_gnd_net_\,
            in3 => \N__26263\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26264\,
            in1 => \_gnd_net_\,
            in2 => \N__15871\,
            in3 => \N__20628\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i3_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20629\,
            in1 => \N__18597\,
            in2 => \_gnd_net_\,
            in3 => \N__26265\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i4_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26266\,
            in1 => \_gnd_net_\,
            in2 => \N__18604\,
            in3 => \N__18627\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i5_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18628\,
            in1 => \N__15840\,
            in2 => \_gnd_net_\,
            in3 => \N__26267\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i6_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26268\,
            in1 => \_gnd_net_\,
            in2 => \N__15847\,
            in3 => \N__15816\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i7_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15817\,
            in1 => \N__15793\,
            in2 => \_gnd_net_\,
            in3 => \N__26269\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => \N__36668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i2_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18767\,
            in1 => \N__22931\,
            in2 => \_gnd_net_\,
            in3 => \N__21040\,
            lcout => \Inst_core.Inst_sync.filteredInput_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37501\,
            ce => 'H',
            sr => \N__18716\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i8_3_lut_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19774\,
            in1 => \N__19756\,
            in2 => \_gnd_net_\,
            in3 => \N__19704\,
            lcout => \GENERIC_FIFO_1.n71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i9_3_lut_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19588\,
            in1 => \N__19564\,
            in2 => \_gnd_net_\,
            in3 => \N__19705\,
            lcout => \GENERIC_FIFO_1.n70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i12_3_lut_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__17983\,
            in1 => \N__17884\,
            in2 => \_gnd_net_\,
            in3 => \N__17695\,
            lcout => \Inst_eia232.Inst_receiver.n3557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i13_3_lut_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010011001"
        )
    port map (
            in0 => \N__17984\,
            in1 => \N__17885\,
            in2 => \_gnd_net_\,
            in3 => \N__17696\,
            lcout => \Inst_eia232.Inst_receiver.n4628\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.busy_87_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__16259\,
            in1 => \N__36425\,
            in2 => \_gnd_net_\,
            in3 => \N__16016\,
            lcout => busy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37508\,
            ce => 'H',
            sr => \N__16208\
        );

    \Inst_eia232.Inst_transmitter.i1_2_lut_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16012\,
            in2 => \_gnd_net_\,
            in3 => \N__16206\,
            lcout => \Inst_eia232.Inst_transmitter.n4634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i3103_2_lut_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16013\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36424\,
            lcout => \Inst_eia232.Inst_transmitter.n4246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__16015\,
            in1 => \N__16207\,
            in2 => \_gnd_net_\,
            in3 => \N__16136\,
            lcout => \Inst_eia232.Inst_transmitter.n8527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i361_2_lut_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36423\,
            in2 => \_gnd_net_\,
            in3 => \N__16068\,
            lcout => \Inst_eia232.Inst_transmitter.n971\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.i3553_2_lut_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16014\,
            in2 => \_gnd_net_\,
            in3 => \N__21683\,
            lcout => \Inst_eia232.Inst_transmitter.n4712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i2_3_lut_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19438\,
            in1 => \N__19413\,
            in2 => \_gnd_net_\,
            in3 => \N__19690\,
            lcout => \GENERIC_FIFO_1.n77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i3_3_lut_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19691\,
            in1 => \N__19360\,
            in2 => \_gnd_net_\,
            in3 => \N__19342\,
            lcout => \GENERIC_FIFO_1.n76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i1_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__22548\,
            in1 => \N__18773\,
            in2 => \_gnd_net_\,
            in3 => \N__22456\,
            lcout => \Inst_core.Inst_sync.filteredInput_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37517\,
            ce => 'H',
            sr => \N__19025\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i4_3_lut_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18979\,
            in1 => \N__19000\,
            in2 => \_gnd_net_\,
            in3 => \N__19664\,
            lcout => \GENERIC_FIFO_1.n75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i5_3_lut_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19258\,
            in1 => \N__19282\,
            in2 => \_gnd_net_\,
            in3 => \N__19665\,
            lcout => \GENERIC_FIFO_1.n74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i6_3_lut_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19666\,
            in1 => \_gnd_net_\,
            in2 => \N__19186\,
            in3 => \N__19213\,
            lcout => \GENERIC_FIFO_1.n73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i6_1_lut_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19178\,
            lcout => \GENERIC_FIFO_1.n1420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921_mux_7_i7_3_lut_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19667\,
            in1 => \_gnd_net_\,
            in2 => \N__19117\,
            in3 => \N__19135\,
            lcout => \GENERIC_FIFO_1.n72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i6_4_lut_adj_120_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19182\,
            in1 => \N__18963\,
            in2 => \N__19563\,
            in3 => \N__17056\,
            lcout => OPEN,
            ltout => \GENERIC_FIFO_1.n16_adj_1279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i5619_4_lut_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__19248\,
            in1 => \N__19414\,
            in2 => \N__16352\,
            in3 => \N__16847\,
            lcout => \GENERIC_FIFO_1.n142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i7_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110111100010"
        )
    port map (
            in0 => \N__23037\,
            in1 => \N__20597\,
            in2 => \N__16289\,
            in3 => \N__19040\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37528\,
            ce => 'H',
            sr => \N__18812\
        );

    \GENERIC_FIFO_1.i7_4_lut_adj_121_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19332\,
            in1 => \N__19745\,
            in2 => \N__17172\,
            in3 => \N__19110\,
            lcout => \GENERIC_FIFO_1.n17_adj_1280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i5_1_lut_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19247\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GENERIC_FIFO_1.n1421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i3_1_lut_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19331\,
            lcout => \GENERIC_FIFO_1.n1423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i4_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__21124\,
            in1 => \N__21151\,
            in2 => \_gnd_net_\,
            in3 => \N__19010\,
            lcout => \Inst_core.Inst_sync.filteredInput_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37539\,
            ce => 'H',
            sr => \N__19505\
        );

    \Inst_eia232.Inst_transmitter.i938_2_lut_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16813\,
            in2 => \_gnd_net_\,
            in3 => \N__16721\,
            lcout => \Inst_eia232.Inst_transmitter.n3608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.i1047_1_lut_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16629\,
            lcout => \GENERIC_FIFO_1.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i2_1_lut_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16579\,
            lcout => \GENERIC_FIFO_1.n1379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i3_1_lut_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16530\,
            lcout => \GENERIC_FIFO_1.n1378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i4_1_lut_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16482\,
            lcout => \GENERIC_FIFO_1.n1377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_675_i7_1_lut_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17115\,
            lcout => \GENERIC_FIFO_1.n1374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_2_lut_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17064\,
            in2 => \N__17018\,
            in3 => \N__17009\,
            lcout => \GENERIC_FIFO_1.n1391\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \GENERIC_FIFO_1.n7938\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_3_lut_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19390\,
            in2 => \N__17006\,
            in3 => \N__16997\,
            lcout => \GENERIC_FIFO_1.n1390\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7938\,
            carryout => \GENERIC_FIFO_1.n7939\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_4_lut_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__16994\,
            in1 => \N__19319\,
            in2 => \N__16988\,
            in3 => \N__16961\,
            lcout => \GENERIC_FIFO_1.n8634\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7939\,
            carryout => \GENERIC_FIFO_1.n7940\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_5_lut_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18961\,
            in2 => \N__16958\,
            in3 => \N__16949\,
            lcout => \GENERIC_FIFO_1.n1388\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7940\,
            carryout => \GENERIC_FIFO_1.n7941\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_6_lut_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__16946\,
            in1 => \N__19235\,
            in2 => \N__16940\,
            in3 => \N__16910\,
            lcout => \GENERIC_FIFO_1.n8628\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7941\,
            carryout => \GENERIC_FIFO_1.n7942\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_7_lut_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16907\,
            in2 => \N__19177\,
            in3 => \N__16895\,
            lcout => \GENERIC_FIFO_1.n1386\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7942\,
            carryout => \GENERIC_FIFO_1.n7943\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_8_lut_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__16892\,
            in1 => \N__19098\,
            in2 => \N__16886\,
            in3 => \N__16865\,
            lcout => \GENERIC_FIFO_1.n8632\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7943\,
            carryout => \GENERIC_FIFO_1.n7944\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_8_THRU_CRY_0_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17349\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7944\,
            carryout => \GENERIC_FIFO_1.n7944_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_9_lut_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__17324\,
            in1 => \N__19729\,
            in2 => \N__17318\,
            in3 => \N__17291\,
            lcout => \GENERIC_FIFO_1.n8630\,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \GENERIC_FIFO_1.n7945\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_10_lut_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19539\,
            in2 => \N__17288\,
            in3 => \N__17276\,
            lcout => \GENERIC_FIFO_1.n1383\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7945\,
            carryout => \GENERIC_FIFO_1.n7946\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.add_676_11_lut_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__17273\,
            in1 => \N__17152\,
            in2 => \N__17267\,
            in3 => \N__17240\,
            lcout => \GENERIC_FIFO_1.n8638\,
            ltout => OPEN,
            carryin => \GENERIC_FIFO_1.n7946\,
            carryout => \GENERIC_FIFO_1.n1392\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.n1392_THRU_LUT4_0_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17237\,
            lcout => \GENERIC_FIFO_1.n1392_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i9_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19682\,
            in1 => \N__17201\,
            in2 => \_gnd_net_\,
            in3 => \N__17154\,
            lcout => \GENERIC_FIFO_1.read_pointer_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i10_1_lut_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17153\,
            lcout => \GENERIC_FIFO_1.n1416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_decoder.executePrev_36_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__17657\,
            in1 => \_gnd_net_\,
            in2 => \N__17967\,
            in3 => \N__17858\,
            lcout => \executePrev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7483_2_lut_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17412\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17653\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n8755_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.state_1__bdd_4_lut_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__17942\,
            in1 => \N__17856\,
            in2 => \N__17378\,
            in3 => \N__17533\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n9123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.state_i1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__17860\,
            in1 => \N__17705\,
            in2 => \N__17375\,
            in3 => \N__17366\,
            lcout => \Inst_eia232.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.i5466_2_lut_4_lut_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__17656\,
            in1 => \N__17372\,
            in2 => \N__17965\,
            in3 => \N__17857\,
            lcout => n1917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7487_2_lut_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__17606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17654\,
            lcout => \Inst_eia232.Inst_receiver.n8784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_2_i6_4_lut_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001111"
        )
    port map (
            in0 => \N__17655\,
            in1 => \N__17534\,
            in2 => \N__17966\,
            in3 => \N__17413\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.state_i2_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__17859\,
            in1 => \N__17946\,
            in2 => \N__17360\,
            in3 => \N__17579\,
            lcout => \Inst_eia232.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i21_3_lut_3_lut_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001000100"
        )
    port map (
            in0 => \N__17662\,
            in1 => \N__17842\,
            in2 => \_gnd_net_\,
            in3 => \N__17603\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7647_3_lut_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__17937\,
            in1 => \_gnd_net_\,
            in2 => \N__17357\,
            in3 => \N__17395\,
            lcout => \Inst_eia232.Inst_receiver.n4767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i4338_4_lut_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__20177\,
            in1 => \N__20210\,
            in2 => \N__17676\,
            in3 => \N__17414\,
            lcout => \Inst_eia232.Inst_receiver.n5505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7481_2_lut_3_lut_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__17604\,
            in1 => \_gnd_net_\,
            in2 => \N__17863\,
            in3 => \N__17663\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n8782_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7653_4_lut_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__17396\,
            in1 => \N__18506\,
            in2 => \N__17399\,
            in3 => \N__17936\,
            lcout => \Inst_eia232.Inst_receiver.n3676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i2_3_lut_adj_99_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17841\,
            in1 => \N__17661\,
            in2 => \_gnd_net_\,
            in3 => \N__20176\,
            lcout => \Inst_eia232.Inst_receiver.n6_adj_1267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_0_i3_4_lut_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111100010111"
        )
    port map (
            in0 => \N__17664\,
            in1 => \N__17938\,
            in2 => \N__18488\,
            in3 => \N__17605\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.state_i0_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__17846\,
            in1 => \N__17950\,
            in2 => \N__17387\,
            in3 => \N__17384\,
            lcout => \Inst_eia232.state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.counter_925__i3_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__17772\,
            in1 => \N__17744\,
            in2 => \N__17441\,
            in3 => \N__17796\,
            lcout => \Inst_eia232.Inst_receiver.counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37542\,
            ce => \N__17567\,
            sr => \N__17552\
        );

    \Inst_eia232.Inst_receiver.counter_925__i2_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__17795\,
            in1 => \_gnd_net_\,
            in2 => \N__17747\,
            in3 => \N__17771\,
            lcout => \Inst_eia232.Inst_receiver.counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37542\,
            ce => \N__17567\,
            sr => \N__17552\
        );

    \Inst_eia232.Inst_receiver.counter_925__i1_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17794\,
            lcout => \Inst_eia232.Inst_receiver.counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37542\,
            ce => \N__17567\,
            sr => \N__17552\
        );

    \Inst_eia232.Inst_receiver.counter_925__i4_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17440\,
            in1 => \N__17459\,
            in2 => \_gnd_net_\,
            in3 => \N__17723\,
            lcout => \Inst_eia232.Inst_receiver.counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37542\,
            ce => \N__17567\,
            sr => \N__17552\
        );

    \Inst_eia232.Inst_receiver.i2_3_lut_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__17768\,
            in1 => \N__17740\,
            in2 => \_gnd_net_\,
            in3 => \N__17793\,
            lcout => \Inst_eia232.Inst_receiver.n3504\,
            ltout => \Inst_eia232.Inst_receiver.n3504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i2_3_lut_adj_86_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17457\,
            in2 => \N__17570\,
            in3 => \N__17434\,
            lcout => \Inst_eia232.Inst_receiver.n957\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.counter_925__i0_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_eia232.Inst_receiver.counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37542\,
            ce => \N__17567\,
            sr => \N__17552\
        );

    \Inst_eia232.Inst_receiver.i5570_3_lut_4_lut_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__17540\,
            in1 => \N__17458\,
            in2 => \N__17675\,
            in3 => \N__17435\,
            lcout => \Inst_eia232.Inst_receiver.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_decoder.wrsize_55_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000010"
        )
    port map (
            in0 => \N__17520\,
            in1 => \N__17503\,
            in2 => \N__18323\,
            in3 => \_gnd_net_\,
            lcout => wrsize,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37531\,
            ce => 'H',
            sr => \N__17486\
        );

    \Inst_core.Inst_decoder.wrspeed_54_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18319\,
            in2 => \N__17507\,
            in3 => \N__18016\,
            lcout => \wrDivider\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37531\,
            ce => 'H',
            sr => \N__17486\
        );

    \Inst_core.Inst_sampler.i857_2_lut_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30992\,
            in2 => \_gnd_net_\,
            in3 => \N__31960\,
            lcout => \Inst_core.Inst_sampler.n1700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i11_4_lut_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20269\,
            in1 => \N__19924\,
            in2 => \N__20030\,
            in3 => \N__19975\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.counter_4__I_0_71_i7_2_lut_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17456\,
            in2 => \_gnd_net_\,
            in3 => \N__17439\,
            lcout => OPEN,
            ltout => \Inst_eia232.Inst_receiver.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i3_4_lut_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__17797\,
            in1 => \N__17773\,
            in2 => \N__17801\,
            in3 => \N__17745\,
            lcout => \Inst_eia232.Inst_receiver.nstate_2_N_133_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i12_4_lut_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20251\,
            in1 => \N__19990\,
            in2 => \N__20234\,
            in3 => \N__20284\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i6596_2_lut_3_lut_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17798\,
            in1 => \N__17774\,
            in2 => \_gnd_net_\,
            in3 => \N__17746\,
            lcout => \Inst_eia232.Inst_receiver.n7777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20507\,
            in1 => \N__22865\,
            in2 => \_gnd_net_\,
            in3 => \N__22435\,
            lcout => \Inst_core.Inst_sync.filteredInput_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37520\,
            ce => 'H',
            sr => \N__18935\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_96_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__17694\,
            in1 => \_gnd_net_\,
            in2 => \N__17982\,
            in3 => \N__17882\,
            lcout => \Inst_eia232.Inst_receiver.n3202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i3313_2_lut_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17971\,
            in2 => \_gnd_net_\,
            in3 => \N__17881\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_adj_107_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17693\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18471\,
            lcout => \Inst_eia232.Inst_receiver.n1_adj_1266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i7571_2_lut_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17692\,
            in2 => \_gnd_net_\,
            in3 => \N__17602\,
            lcout => \Inst_eia232.Inst_receiver.n8826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i5549_2_lut_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36658\,
            in2 => \_gnd_net_\,
            in3 => \N__25367\,
            lcout => \Inst_core.n6713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_prescaler.i5470_2_lut_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18568\,
            in2 => \_gnd_net_\,
            in3 => \N__18535\,
            lcout => \Inst_eia232.Inst_prescaler.counter_4__N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_adj_80_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18416\,
            in2 => \_gnd_net_\,
            in3 => \N__18380\,
            lcout => n12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i3_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__18080\,
            in1 => \N__18239\,
            in2 => \N__18202\,
            in3 => \N__34701\,
            lcout => \Inst_eia232.Inst_receiver.cmd_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i2_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__18237\,
            in1 => \N__18303\,
            in2 => \N__18198\,
            in3 => \N__34706\,
            lcout => \Inst_eia232.Inst_receiver.cmd_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.opcode_i1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__18114\,
            in1 => \N__34699\,
            in2 => \N__18318\,
            in3 => \N__18238\,
            lcout => \Inst_eia232.Inst_receiver.cmd_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18173\,
            in1 => \N__18113\,
            in2 => \_gnd_net_\,
            in3 => \N__18079\,
            lcout => \Inst_eia232.Inst_receiver.n69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i27_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__28192\,
            in1 => \N__35633\,
            in2 => \N__35067\,
            in3 => \N__34700\,
            lcout => cmd_34,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_109_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__17975\,
            in1 => \N__20091\,
            in2 => \_gnd_net_\,
            in3 => \N__17883\,
            lcout => \Inst_eia232.Inst_receiver.n8376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i5_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29097\,
            in1 => \N__34698\,
            in2 => \N__31397\,
            in3 => \N__35059\,
            lcout => cmd_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_prescaler.scaled_28_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18572\,
            in2 => \_gnd_net_\,
            in3 => \N__18539\,
            lcout => \trxClock\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i3_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26712\,
            in1 => \N__20689\,
            in2 => \_gnd_net_\,
            in3 => \N__18640\,
            lcout => \valueRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i3_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21865\,
            in1 => \N__26711\,
            in2 => \_gnd_net_\,
            in3 => \N__18895\,
            lcout => \maskRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i22_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29757\,
            in1 => \N__35790\,
            in2 => \_gnd_net_\,
            in3 => \N__18735\,
            lcout => \configRegister_23_adj_1339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i22_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26026\,
            in1 => \N__29758\,
            in2 => \_gnd_net_\,
            in3 => \N__18659\,
            lcout => \configRegister_23_adj_1379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i2_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__34817\,
            in1 => \N__29706\,
            in2 => \N__34205\,
            in3 => \N__34996\,
            lcout => cmd_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i32_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__34995\,
            in1 => \N__20446\,
            in2 => \N__18470\,
            in3 => \N__34818\,
            lcout => cmd_39,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_7706_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__21818\,
            in1 => \N__23026\,
            in2 => \N__30467\,
            in3 => \N__20410\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_bdd_4_lut_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__20412\,
            in1 => \N__28081\,
            in2 => \N__18437\,
            in3 => \N__25490\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9096_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_754_i1_3_lut_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__21932\,
            in1 => \N__21466\,
            in2 => \N__18665\,
            in3 => \N__18658\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__32343\,
            in1 => \N__30923\,
            in2 => \N__20414\,
            in3 => \N__21817\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_bdd_4_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__33646\,
            in1 => \N__31794\,
            in2 => \N__18662\,
            in3 => \N__20411\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_746_i1_3_lut_4_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__18657\,
            in1 => \N__21931\,
            in2 => \N__18644\,
            in3 => \N__21487\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i3_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110010101101010"
        )
    port map (
            in0 => \N__18641\,
            in1 => \N__18629\,
            in2 => \N__20593\,
            in3 => \N__32344\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37488\,
            ce => 'H',
            sr => \N__18881\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i2_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110111100010"
        )
    port map (
            in0 => \N__30922\,
            in1 => \N__20576\,
            in2 => \N__18605\,
            in3 => \N__18707\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37504\,
            ce => 'H',
            sr => \N__18911\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_7697_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__20482\,
            in1 => \N__32338\,
            in2 => \N__21959\,
            in3 => \N__30921\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_bdd_4_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__31789\,
            in1 => \N__33634\,
            in2 => \N__18578\,
            in3 => \N__21957\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9084_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_730_i1_3_lut_4_lut_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__18736\,
            in1 => \N__22108\,
            in2 => \N__18575\,
            in3 => \N__24973\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelL16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__23025\,
            in1 => \N__20483\,
            in2 => \N__30466\,
            in3 => \N__21956\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_bdd_4_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__21958\,
            in1 => \N__28077\,
            in2 => \N__18740\,
            in3 => \N__25489\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n9090_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_738_i1_3_lut_4_lut_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__22109\,
            in1 => \N__18737\,
            in2 => \N__18719\,
            in3 => \N__24928\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.i3571_1_lut_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21014\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22025\,
            in1 => \N__35988\,
            in2 => \_gnd_net_\,
            in3 => \N__18800\,
            lcout => \maskRegister_0_adj_1288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20699\,
            in1 => \N__29714\,
            in2 => \_gnd_net_\,
            in3 => \N__18706\,
            lcout => \valueRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i23_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22226\,
            in1 => \N__29290\,
            in2 => \_gnd_net_\,
            in3 => \N__20845\,
            lcout => \configRegister_24_adj_1298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i24_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35643\,
            in1 => \_gnd_net_\,
            in2 => \N__34098\,
            in3 => \N__20554\,
            lcout => \configRegister_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i5_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18691\,
            in1 => \N__20700\,
            in2 => \_gnd_net_\,
            in3 => \N__31369\,
            lcout => \valueRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i23_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34046\,
            in1 => \N__18676\,
            in2 => \_gnd_net_\,
            in3 => \N__22225\,
            lcout => \configRegister_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3483_1_lut_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18799\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i7_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18824\,
            in1 => \N__27201\,
            in2 => \_gnd_net_\,
            in3 => \N__21887\,
            lcout => \maskRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22558\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i6_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34408\,
            in1 => \N__21886\,
            in2 => \_gnd_net_\,
            in3 => \N__18848\,
            lcout => \maskRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i2_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22930\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i6_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34409\,
            in1 => \N__20695\,
            in2 => \_gnd_net_\,
            in3 => \N__18751\,
            lcout => \valueRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i7_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27200\,
            in1 => \_gnd_net_\,
            in2 => \N__34501\,
            in3 => \N__23089\,
            lcout => \valueRegister_7_adj_1289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i2_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29707\,
            in1 => \N__21884\,
            in2 => \_gnd_net_\,
            in3 => \N__18923\,
            lcout => \maskRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i4_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21885\,
            in1 => \N__29110\,
            in2 => \_gnd_net_\,
            in3 => \N__18872\,
            lcout => \maskRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__19514\,
            in1 => \N__22318\,
            in2 => \_gnd_net_\,
            in3 => \N__22636\,
            lcout => \Inst_core.Inst_sync.filteredInput_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37530\,
            ce => 'H',
            sr => \N__20969\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3581_1_lut_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18922\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4740\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3582_1_lut_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18896\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3583_1_lut_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18871\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4742\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3585_1_lut_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18847\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3586_1_lut_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18823\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_1_lut_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36812\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.n3670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i1_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23302\,
            lcout => \Inst_core.Inst_sync.demuxedInput_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i7_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27206\,
            in1 => \N__22027\,
            in2 => \_gnd_net_\,
            in3 => \N__26932\,
            lcout => \maskRegister_7_adj_1281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i4_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20691\,
            in1 => \N__19060\,
            in2 => \_gnd_net_\,
            in3 => \N__29115\,
            lcout => \valueRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i7_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27205\,
            in1 => \N__31111\,
            in2 => \_gnd_net_\,
            in3 => \N__24867\,
            lcout => divider_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i7_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31110\,
            in1 => \N__23018\,
            in2 => \N__22493\,
            in3 => \N__31964\,
            lcout => \memoryOut_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i2_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22026\,
            in1 => \N__29679\,
            in2 => \_gnd_net_\,
            in3 => \N__20909\,
            lcout => \maskRegister_2_adj_1286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i4_1_lut_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18962\,
            lcout => \GENERIC_FIFO_1.n1422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i7_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19036\,
            in1 => \N__27209\,
            in2 => \_gnd_net_\,
            in3 => \N__20701\,
            lcout => \valueRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.i3570_1_lut_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22895\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i4_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21152\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i3_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19004\,
            in1 => \N__18969\,
            in2 => \_gnd_net_\,
            in3 => \N__19700\,
            lcout => \GENERIC_FIFO_1.read_pointer_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.i3572_1_lut_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i2_1_lut_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19391\,
            lcout => \GENERIC_FIFO_1.n1424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i7_1_lut_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19099\,
            lcout => \GENERIC_FIFO_1.n1419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i1_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19442\,
            in1 => \N__19400\,
            in2 => \_gnd_net_\,
            in3 => \N__19683\,
            lcout => \GENERIC_FIFO_1.read_pointer_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i2_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19684\,
            in1 => \N__19364\,
            in2 => \_gnd_net_\,
            in3 => \N__19330\,
            lcout => \GENERIC_FIFO_1.read_pointer_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.inv_692_i9_1_lut_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19540\,
            lcout => \GENERIC_FIFO_1.n1417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i4_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19685\,
            in1 => \N__19286\,
            in2 => \_gnd_net_\,
            in3 => \N__19246\,
            lcout => \GENERIC_FIFO_1.read_pointer_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i5_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19217\,
            in1 => \N__19176\,
            in2 => \_gnd_net_\,
            in3 => \N__19686\,
            lcout => \GENERIC_FIFO_1.read_pointer_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i6_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19687\,
            in1 => \N__19139\,
            in2 => \_gnd_net_\,
            in3 => \N__19109\,
            lcout => \GENERIC_FIFO_1.read_pointer_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i7_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19781\,
            in1 => \N__19741\,
            in2 => \_gnd_net_\,
            in3 => \N__19688\,
            lcout => \GENERIC_FIFO_1.read_pointer_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GENERIC_FIFO_1.read_pointer_921__i8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19689\,
            in1 => \_gnd_net_\,
            in2 => \N__19553\,
            in3 => \N__19592\,
            lcout => \GENERIC_FIFO_1.read_pointer_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i0_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22317\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.i3573_1_lut_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19493\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4732\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input180Delay_i5_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23126\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input180Delay_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input180Delay_i6_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23165\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input180Delay_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i4_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21263\,
            lcout => \Inst_core.Inst_sync.synchronizedInput_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input180Delay_i4_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21241\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input180Delay_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i0_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22685\,
            lcout => \Inst_core.Inst_sync.demuxedInput_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i1_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19480\,
            in2 => \_gnd_net_\,
            in3 => \N__19469\,
            lcout => testcnt_c_0,
            ltout => OPEN,
            carryin => \bfn_6_1_0_\,
            carryout => n7862,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i2_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19903\,
            in2 => \_gnd_net_\,
            in3 => \N__19892\,
            lcout => testcnt_c_1,
            ltout => OPEN,
            carryin => n7862,
            carryout => n7863,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i3_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19882\,
            in2 => \_gnd_net_\,
            in3 => \N__19871\,
            lcout => testcnt_c_2,
            ltout => OPEN,
            carryin => n7863,
            carryout => n7864,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i4_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19867\,
            in2 => \_gnd_net_\,
            in3 => \N__19856\,
            lcout => testcnt_c_3,
            ltout => OPEN,
            carryin => n7864,
            carryout => n7865,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i5_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19852\,
            in2 => \_gnd_net_\,
            in3 => \N__19841\,
            lcout => testcnt_c_4,
            ltout => OPEN,
            carryin => n7865,
            carryout => n7866,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i6_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19837\,
            in2 => \_gnd_net_\,
            in3 => \N__19826\,
            lcout => testcnt_c_5,
            ltout => OPEN,
            carryin => n7866,
            carryout => n7867,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i7_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19816\,
            in2 => \_gnd_net_\,
            in3 => \N__19805\,
            lcout => testcnt_c_6,
            ltout => OPEN,
            carryin => n7867,
            carryout => n7868,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testcnt_i_917__i8_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19792\,
            in2 => \_gnd_net_\,
            in3 => \N__19802\,
            lcout => testcnt_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i9_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20011\,
            in1 => \N__26114\,
            in2 => \_gnd_net_\,
            in3 => \N__23998\,
            lcout => \configRegister_8_adj_1392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i2_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26113\,
            in1 => \N__19957\,
            in2 => \_gnd_net_\,
            in3 => \N__34267\,
            lcout => \configRegister_1_adj_1399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i3_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29625\,
            in1 => \N__19939\,
            in2 => \_gnd_net_\,
            in3 => \N__26118\,
            lcout => \configRegister_2_adj_1398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i2_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35800\,
            in1 => \N__23374\,
            in2 => \_gnd_net_\,
            in3 => \N__34266\,
            lcout => \configRegister_1_adj_1359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i3_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29624\,
            in1 => \N__23344\,
            in2 => \_gnd_net_\,
            in3 => \N__35801\,
            lcout => \configRegister_2_adj_1358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i4_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26721\,
            in1 => \_gnd_net_\,
            in2 => \N__26134\,
            in3 => \N__20053\,
            lcout => \configRegister_3_adj_1397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i4_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35802\,
            in1 => \N__23314\,
            in2 => \_gnd_net_\,
            in3 => \N__26720\,
            lcout => \configRegister_3_adj_1357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i3_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29623\,
            in1 => \N__34776\,
            in2 => \N__26732\,
            in3 => \N__35045\,
            lcout => cmd_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20498\,
            in1 => \N__25082\,
            in2 => \N__21404\,
            in3 => \N__19961\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7914\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i1_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__19958\,
            in1 => \N__21437\,
            in2 => \N__25321\,
            in3 => \N__19946\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7914\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7915\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i2_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__19943\,
            in1 => \N__25293\,
            in2 => \N__19928\,
            in3 => \N__19913\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7915\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7916\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i3_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20054\,
            in1 => \N__21347\,
            in2 => \N__25322\,
            in3 => \N__20042\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7916\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7917\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i4_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__20465\,
            in1 => \N__25297\,
            in2 => \N__21424\,
            in3 => \N__20039\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7917\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7918\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i5_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21287\,
            in1 => \N__21334\,
            in2 => \N__25323\,
            in3 => \N__20036\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7918\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7919\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i6_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__20354\,
            in1 => \N__25301\,
            in2 => \N__21452\,
            in3 => \N__20033\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7919\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7920\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i7_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20324\,
            in1 => \N__20029\,
            in2 => \N__25324\,
            in3 => \N__20015\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7920\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7921\,
            clk => \N__37556\,
            ce => \N__25697\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i8_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20012\,
            in1 => \N__21320\,
            in2 => \N__25325\,
            in3 => \N__19997\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7922\,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i9_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__24083\,
            in1 => \N__25308\,
            in2 => \N__19994\,
            in3 => \N__19979\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7922\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7923\,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i10_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21506\,
            in1 => \N__19976\,
            in2 => \N__25326\,
            in3 => \N__19964\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7923\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7924\,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i11_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__21518\,
            in1 => \N__25312\,
            in2 => \N__20288\,
            in3 => \N__20273\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7924\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7925\,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i12_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23882\,
            in1 => \N__20270\,
            in2 => \N__25327\,
            in3 => \N__20258\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7925\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7926\,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i13_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__26162\,
            in1 => \N__25316\,
            in2 => \N__21362\,
            in3 => \N__20255\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7926\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7927\,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i14_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__25547\,
            in1 => \N__20252\,
            in2 => \N__25328\,
            in3 => \N__20240\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7927\,
            carryout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7928\,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i15_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__20233\,
            in1 => \N__25320\,
            in2 => \N__21773\,
            in3 => \N__20237\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37544\,
            ce => \N__25696\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.bytecount_i0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__20115\,
            in1 => \N__20219\,
            in2 => \_gnd_net_\,
            in3 => \N__20186\,
            lcout => \Inst_eia232.Inst_receiver.bytecount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37533\,
            ce => \N__20099\,
            sr => \N__20060\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3603_1_lut_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20335\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3604_1_lut_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3606_1_lut_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20389\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3607_1_lut_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20377\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i6_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34404\,
            in2 => \N__23921\,
            in3 => \N__20390\,
            lcout => \maskRegister_6_adj_1362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i7_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20378\,
            in1 => \N__27141\,
            in2 => \_gnd_net_\,
            in3 => \N__23916\,
            lcout => \maskRegister_7_adj_1361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i4_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23912\,
            in1 => \N__29063\,
            in2 => \_gnd_net_\,
            in3 => \N__20366\,
            lcout => \maskRegister_4_adj_1364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i7_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__26048\,
            in1 => \N__20347\,
            in2 => \N__34429\,
            in3 => \_gnd_net_\,
            lcout => \configRegister_6_adj_1394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i3_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23911\,
            in1 => \N__26653\,
            in2 => \_gnd_net_\,
            in3 => \N__20336\,
            lcout => \maskRegister_3_adj_1365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i8_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26049\,
            in1 => \N__20320\,
            in2 => \_gnd_net_\,
            in3 => \N__27142\,
            lcout => \configRegister_7_adj_1393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__27140\,
            in1 => \N__34702\,
            in2 => \N__23992\,
            in3 => \N__35058\,
            lcout => cmd_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i9_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__35057\,
            in1 => \N__23974\,
            in2 => \N__34777\,
            in3 => \N__26596\,
            lcout => cmd_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34522\,
            in1 => \N__35926\,
            in2 => \_gnd_net_\,
            in3 => \N__20299\,
            lcout => \valueRegister_0_adj_1296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i3_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22864\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i21_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29331\,
            in1 => \N__24179\,
            in2 => \_gnd_net_\,
            in3 => \N__20721\,
            lcout => \configRegister_22_adj_1300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i1_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21888\,
            in1 => \N__34179\,
            in2 => \_gnd_net_\,
            in3 => \N__20956\,
            lcout => \maskRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i1_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26100\,
            in1 => \N__35927\,
            in2 => \_gnd_net_\,
            in3 => \N__20497\,
            lcout => \configRegister_0_adj_1400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i19_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35794\,
            in1 => \N__26535\,
            in2 => \_gnd_net_\,
            in3 => \N__20481\,
            lcout => \configRegister_20_adj_1342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i5_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26101\,
            in1 => \N__20461\,
            in2 => \_gnd_net_\,
            in3 => \N__29064\,
            lcout => \configRegister_4_adj_1396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i15_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35364\,
            in1 => \N__20445\,
            in2 => \_gnd_net_\,
            in3 => \N__22378\,
            lcout => fwd_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3482_1_lut_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21829\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i20_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24664\,
            in1 => \N__26119\,
            in2 => \_gnd_net_\,
            in3 => \N__20413\,
            lcout => \configRegister_21_adj_1381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i22_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29300\,
            in1 => \N__29751\,
            in2 => \_gnd_net_\,
            in3 => \N__20738\,
            lcout => \configRegister_23_adj_1299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22037\,
            in1 => \N__26716\,
            in2 => \_gnd_net_\,
            in3 => \N__20896\,
            lcout => \maskRegister_3_adj_1285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i20_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29299\,
            in1 => \N__24663\,
            in2 => \_gnd_net_\,
            in3 => \N__20763\,
            lcout => \configRegister_21_adj_1301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i22_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24662\,
            in1 => \N__34775\,
            in2 => \N__24178\,
            in3 => \N__34965\,
            lcout => cmd_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i5_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34523\,
            in1 => \N__24328\,
            in2 => \_gnd_net_\,
            in3 => \N__31387\,
            lcout => \valueRegister_5_adj_1291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20702\,
            in1 => \N__34196\,
            in2 => \_gnd_net_\,
            in3 => \N__20615\,
            lcout => \valueRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_722_i1_3_lut_4_lut_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__20737\,
            in1 => \N__20774\,
            in2 => \N__20819\,
            in3 => \N__20723\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000111100"
        )
    port map (
            in0 => \N__20633\,
            in1 => \N__20614\,
            in2 => \N__33652\,
            in3 => \N__20561\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37513\,
            ce => 'H',
            sr => \N__20942\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__23039\,
            in1 => \N__20863\,
            in2 => \N__20765\,
            in3 => \N__30456\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_bdd_4_lut_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__25488\,
            in1 => \N__28028\,
            in2 => \N__20777\,
            in3 => \N__20762\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9078\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_7688_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__30924\,
            in1 => \N__32339\,
            in2 => \N__20764\,
            in3 => \N__20862\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_bdd_4_lut_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__31790\,
            in1 => \N__33638\,
            in2 => \N__20768\,
            in3 => \N__20761\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_714_i1_3_lut_4_lut_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__20736\,
            in1 => \N__20722\,
            in2 => \N__20705\,
            in3 => \N__20833\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_flags.filter_16_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34226\,
            in1 => \N__22260\,
            in2 => \_gnd_net_\,
            in3 => \N__22583\,
            lcout => \flagFilter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i5_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22035\,
            in1 => \N__31368\,
            in2 => \_gnd_net_\,
            in3 => \N__20878\,
            lcout => \maskRegister_5_adj_1283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i4_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__35365\,
            in1 => \N__26519\,
            in2 => \N__24239\,
            in3 => \_gnd_net_\,
            lcout => fwd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29109\,
            in1 => \N__34529\,
            in2 => \_gnd_net_\,
            in3 => \N__24550\,
            lcout => \valueRegister_4_adj_1292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i1_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34227\,
            in1 => \N__22034\,
            in2 => \_gnd_net_\,
            in3 => \N__20923\,
            lcout => \maskRegister_1_adj_1287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i21_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__26518\,
            in1 => \N__34841\,
            in2 => \N__24684\,
            in3 => \N__35056\,
            lcout => cmd_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i23_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35832\,
            in1 => \N__24949\,
            in2 => \_gnd_net_\,
            in3 => \N__22218\,
            lcout => \configRegister_24_adj_1338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i19_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26520\,
            in1 => \N__29326\,
            in2 => \_gnd_net_\,
            in3 => \N__20864\,
            lcout => \configRegister_20_adj_1302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__26356\,
            in1 => \N__20818\,
            in2 => \N__20849\,
            in3 => \N__20834\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20817\,
            in1 => \N__20790\,
            in2 => \_gnd_net_\,
            in3 => \N__26349\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26350\,
            in1 => \_gnd_net_\,
            in2 => \N__20797\,
            in3 => \N__22122\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i3_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22123\,
            in1 => \N__29802\,
            in2 => \_gnd_net_\,
            in3 => \N__26351\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i4_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26352\,
            in1 => \_gnd_net_\,
            in2 => \N__29809\,
            in3 => \N__26856\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i5_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26857\,
            in1 => \N__24573\,
            in2 => \_gnd_net_\,
            in3 => \N__26353\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i6_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26354\,
            in1 => \_gnd_net_\,
            in2 => \N__24580\,
            in3 => \N__24309\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i7_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24310\,
            in1 => \N__30244\,
            in2 => \_gnd_net_\,
            in3 => \N__26355\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => \N__36609\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i6_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20995\,
            in1 => \N__22514\,
            in2 => \_gnd_net_\,
            in3 => \N__22712\,
            lcout => \Inst_core.Inst_sync.filteredInput_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37543\,
            ce => 'H',
            sr => \N__21080\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3587_1_lut_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20924\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4746\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3588_1_lut_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20908\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3589_1_lut_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20897\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3590_1_lut_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20980\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3591_1_lut_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20882\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4750\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_demux.output_6__12_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.demuxedInput_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i4_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29107\,
            in2 => \N__31136\,
            in3 => \N__27360\,
            lcout => divider_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i2_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31106\,
            in1 => \N__30909\,
            in2 => \N__21023\,
            in3 => \N__31963\,
            lcout => \memoryOut_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.i1680_3_lut_4_lut_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__23239\,
            in1 => \N__22596\,
            in2 => \N__21047\,
            in3 => \N__26380\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sync.n2789_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i2_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22920\,
            in1 => \_gnd_net_\,
            in2 => \N__21026\,
            in3 => \N__22804\,
            lcout => \syncedInput_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i6_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__22721\,
            in1 => \N__21010\,
            in2 => \N__20996\,
            in3 => \N__22750\,
            lcout => \syncedInput_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i4_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29108\,
            in1 => \N__22036\,
            in2 => \_gnd_net_\,
            in3 => \N__20981\,
            lcout => \maskRegister_4_adj_1284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i5_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__21178\,
            in1 => \N__22529\,
            in2 => \_gnd_net_\,
            in3 => \N__22827\,
            lcout => \Inst_core.Inst_sync.filteredInput_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37569\,
            ce => 'H',
            sr => \N__21059\
        );

    \Inst_core.Inst_sync.Inst_filter.i3478_1_lut_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21109\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.i3576_1_lut_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20930\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i3580_1_lut_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20957\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input180Delay_i7_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23111\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input180Delay_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i4_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31104\,
            in1 => \N__28027\,
            in2 => \N__21095\,
            in3 => \N__31961\,
            lcout => \memoryOut_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_demux.output_4__14_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22660\,
            lcout => \Inst_core.Inst_sync.demuxedInput_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.n2566_bdd_4_lut_7720_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__22807\,
            in1 => \N__22764\,
            in2 => \N__22832\,
            in3 => \N__23122\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sync.n9063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i5_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__22766\,
            in1 => \N__21179\,
            in2 => \N__21164\,
            in3 => \N__22894\,
            lcout => \syncedInput_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i5_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31105\,
            in1 => \N__25455\,
            in2 => \N__21161\,
            in3 => \N__31962\,
            lcout => \memoryOut_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.n2566_bdd_4_lut_7679_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__22763\,
            in1 => \N__21144\,
            in2 => \N__21242\,
            in3 => \N__22808\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sync.n9057_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i4_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__21131\,
            in1 => \N__21110\,
            in2 => \N__21098\,
            in3 => \N__22765\,
            lcout => \syncedInput_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.i3575_1_lut_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21086\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.i3574_1_lut_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21065\,
            lcout => \Inst_core.Inst_sync.Inst_filter.n4733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i4_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21259\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.match_84_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23642\,
            lcout => \Inst_core.Inst_trigger.stageMatch_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37596\,
            ce => \N__32609\,
            sr => \N__23411\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i6_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__21800\,
            in1 => \N__21302\,
            in2 => \N__33557\,
            in3 => \N__30457\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37585\,
            ce => 'H',
            sr => \N__21227\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i9_4_lut_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23527\,
            in1 => \N__23362\,
            in2 => \N__23573\,
            in3 => \N__23392\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i15_4_lut_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21185\,
            in1 => \N__21206\,
            in2 => \N__21215\,
            in3 => \N__21212\,
            lcout => \Inst_core.n31_adj_1174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i11_4_lut_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23332\,
            in1 => \N__23821\,
            in2 => \N__23512\,
            in3 => \N__23446\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i10_4_lut_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23803\,
            in1 => \N__23587\,
            in2 => \N__23552\,
            in3 => \N__23491\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i7_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100101101100"
        )
    port map (
            in0 => \N__33538\,
            in1 => \N__21275\,
            in2 => \N__21785\,
            in3 => \N__23053\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37572\,
            ce => 'H',
            sr => \N__21200\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i12_4_lut_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23788\,
            in1 => \N__23473\,
            in2 => \N__23684\,
            in3 => \N__23428\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i9_4_lut_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21448\,
            in1 => \N__21436\,
            in2 => \N__21425\,
            in3 => \N__21400\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i15_4_lut_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21389\,
            in1 => \N__21308\,
            in2 => \N__21377\,
            in3 => \N__21374\,
            lcout => \Inst_core.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i10_4_lut_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21358\,
            in1 => \N__21346\,
            in2 => \N__21335\,
            in3 => \N__21319\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i6_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36088\,
            in1 => \N__34424\,
            in2 => \_gnd_net_\,
            in3 => \N__21298\,
            lcout => \valueRegister_6_adj_1370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i12_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34593\,
            in1 => \N__29267\,
            in2 => \_gnd_net_\,
            in3 => \N__28405\,
            lcout => \configRegister_11_adj_1309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i6_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31402\,
            in1 => \N__21286\,
            in2 => \_gnd_net_\,
            in3 => \N__26088\,
            lcout => \configRegister_5_adj_1395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i11_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35799\,
            in1 => \N__25588\,
            in2 => \_gnd_net_\,
            in3 => \N__23458\,
            lcout => \configRegister_10_adj_1350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i11_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__25587\,
            in1 => \N__34594\,
            in2 => \N__34840\,
            in3 => \N__35068\,
            lcout => cmd_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i7_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36089\,
            in1 => \N__27198\,
            in2 => \_gnd_net_\,
            in3 => \N__21274\,
            lcout => \valueRegister_7_adj_1369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i12_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34595\,
            in1 => \N__26087\,
            in2 => \_gnd_net_\,
            in3 => \N__21517\,
            lcout => \configRegister_11_adj_1389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i11_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26086\,
            in1 => \N__25589\,
            in2 => \_gnd_net_\,
            in3 => \N__21505\,
            lcout => \configRegister_10_adj_1390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__26342\,
            in1 => \N__21473\,
            in2 => \N__21494\,
            in3 => \N__21755\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i1_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21472\,
            in1 => \N__31701\,
            in2 => \_gnd_net_\,
            in3 => \N__26335\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i2_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__26336\,
            in1 => \N__33456\,
            in2 => \N__31708\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33457\,
            in1 => \N__28635\,
            in2 => \_gnd_net_\,
            in3 => \N__26337\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i4_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26338\,
            in1 => \_gnd_net_\,
            in2 => \N__28642\,
            in3 => \N__32373\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i5_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32374\,
            in1 => \N__28113\,
            in2 => \_gnd_net_\,
            in3 => \N__26339\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i6_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26340\,
            in1 => \_gnd_net_\,
            in2 => \N__28120\,
            in3 => \N__25527\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i7_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25528\,
            in1 => \N__21796\,
            in2 => \_gnd_net_\,
            in3 => \N__26341\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => \N__36643\,
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i4_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__35060\,
            in1 => \N__26652\,
            in2 => \N__29128\,
            in3 => \N__34796\,
            lcout => cmd_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i16_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33913\,
            in1 => \N__26076\,
            in2 => \_gnd_net_\,
            in3 => \N__21766\,
            lcout => \configRegister_15_adj_1385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i9_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__23978\,
            in1 => \_gnd_net_\,
            in2 => \N__28489\,
            in3 => \N__29333\,
            lcout => \configRegister_8_adj_1312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i23_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26075\,
            in1 => \N__21754\,
            in2 => \_gnd_net_\,
            in3 => \N__22219\,
            lcout => \configRegister_24_adj_1378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i5_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23917\,
            in1 => \N__31352\,
            in2 => \_gnd_net_\,
            in3 => \N__25639\,
            lcout => \maskRegister_5_adj_1363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.disabledGroupsReg_i0_i0_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22285\,
            in1 => \N__29676\,
            in2 => \_gnd_net_\,
            in3 => \N__21547\,
            lcout => \disabledGroupsReg_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_transmitter.disabledBuffer_i0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__21731\,
            in1 => \N__21681\,
            in2 => \N__21551\,
            in3 => \N__21532\,
            lcout => \Inst_eia232.Inst_transmitter.disabledBuffer_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i24_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__35050\,
            in1 => \N__22203\,
            in2 => \N__29756\,
            in3 => \N__34801\,
            lcout => cmd_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__34206\,
            in1 => \N__34800\,
            in2 => \N__35954\,
            in3 => \N__35051\,
            lcout => cmd_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i14_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29383\,
            in1 => \N__34106\,
            in2 => \_gnd_net_\,
            in3 => \N__33835\,
            lcout => \configRegister_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i6_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29457\,
            in1 => \N__34410\,
            in2 => \_gnd_net_\,
            in3 => \N__27394\,
            lcout => \valueRegister_6_adj_1330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i14_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29384\,
            in1 => \N__29332\,
            in2 => \_gnd_net_\,
            in3 => \N__28804\,
            lcout => \configRegister_13_adj_1307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i21_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24175\,
            in1 => \N__26102\,
            in2 => \_gnd_net_\,
            in3 => \N__21925\,
            lcout => \configRegister_22_adj_1380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i22_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29745\,
            in1 => \N__34107\,
            in2 => \_gnd_net_\,
            in3 => \N__21904\,
            lcout => \configRegister_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i8_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31197\,
            in1 => \N__23985\,
            in2 => \_gnd_net_\,
            in3 => \N__27262\,
            lcout => divider_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i8_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35476\,
            in1 => \N__23997\,
            in2 => \_gnd_net_\,
            in3 => \N__24265\,
            lcout => bwd_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21890\,
            in1 => \N__35925\,
            in2 => \_gnd_net_\,
            in3 => \N__21830\,
            lcout => \maskRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i19_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26112\,
            in1 => \N__26536\,
            in2 => \_gnd_net_\,
            in3 => \N__21816\,
            lcout => \configRegister_20_adj_1382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i21_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24153\,
            in1 => \N__35795\,
            in2 => \_gnd_net_\,
            in3 => \N__22102\,
            lcout => \configRegister_22_adj_1340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i25_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__34797\,
            in1 => \N__24101\,
            in2 => \N__22216\,
            in3 => \N__34959\,
            lcout => cmd_32,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i30_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__34958\,
            in1 => \N__24061\,
            in2 => \N__24390\,
            in3 => \N__34798\,
            lcout => cmd_37,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i11_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34582\,
            in1 => \N__31196\,
            in2 => \_gnd_net_\,
            in3 => \N__30771\,
            lcout => divider_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i20_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22061\,
            in1 => \N__24668\,
            in2 => \_gnd_net_\,
            in3 => \N__34084\,
            lcout => \configRegister_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i6_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22024\,
            in1 => \N__34422\,
            in2 => \_gnd_net_\,
            in3 => \N__29779\,
            lcout => \maskRegister_6_adj_1282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34527\,
            in1 => \N__34231\,
            in2 => \_gnd_net_\,
            in3 => \N__22135\,
            lcout => \valueRegister_1_adj_1295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i9_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26586\,
            in1 => \N__31185\,
            in2 => \_gnd_net_\,
            in3 => \N__24888\,
            lcout => divider_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i20_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35820\,
            in1 => \N__24669\,
            in2 => \_gnd_net_\,
            in3 => \N__21952\,
            lcout => \configRegister_21_adj_1341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i16_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__35017\,
            in1 => \N__33898\,
            in2 => \N__36184\,
            in3 => \N__34804\,
            lcout => cmd_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_flags.inverted_18_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22615\,
            in1 => \N__27191\,
            in2 => \_gnd_net_\,
            in3 => \N__22278\,
            lcout => \flagInverted\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i8_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22217\,
            in1 => \N__35406\,
            in2 => \_gnd_net_\,
            in3 => \N__24436\,
            lcout => fwd_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i11_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28177\,
            in1 => \_gnd_net_\,
            in2 => \N__35441\,
            in3 => \N__24251\,
            lcout => fwd_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i5_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35407\,
            in1 => \N__24685\,
            in2 => \_gnd_net_\,
            in3 => \N__22346\,
            lcout => fwd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i20_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31164\,
            in1 => \_gnd_net_\,
            in2 => \N__26534\,
            in3 => \N__25050\,
            lcout => divider_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i5_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31351\,
            in1 => \N__35401\,
            in2 => \_gnd_net_\,
            in3 => \N__26785\,
            lcout => bwd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i6_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35405\,
            in1 => \N__24176\,
            in2 => \_gnd_net_\,
            in3 => \N__22361\,
            lcout => fwd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i22_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24177\,
            in1 => \N__31165\,
            in2 => \_gnd_net_\,
            in3 => \N__32046\,
            lcout => divider_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i19_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26524\,
            in1 => \N__34120\,
            in2 => \_gnd_net_\,
            in3 => \N__22161\,
            lcout => \configRegister_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i1_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001011010"
        )
    port map (
            in0 => \N__22142\,
            in1 => \N__22124\,
            in2 => \N__33645\,
            in3 => \N__30359\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37545\,
            ce => 'H',
            sr => \N__22400\
        );

    \Inst_core.Inst_controller.i10_4_lut_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24449\,
            in1 => \N__24185\,
            in2 => \N__30173\,
            in3 => \N__24470\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_controller.n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i1_4_lut_adj_55_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__37663\,
            in1 => \N__22382\,
            in2 => \N__22364\,
            in3 => \N__24218\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_controller.n4_adj_986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i1_4_lut_adj_56_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__22360\,
            in1 => \N__36989\,
            in2 => \N__22349\,
            in3 => \N__22331\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_controller.n4_adj_987_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i1_4_lut_adj_57_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111111"
        )
    port map (
            in0 => \N__37025\,
            in1 => \N__22345\,
            in2 => \N__22334\,
            in3 => \N__29861\,
            lcout => \Inst_core.Inst_controller.nstate_1_N_829_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i15_2_lut_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24035\,
            in2 => \_gnd_net_\,
            in3 => \N__37697\,
            lcout => \Inst_core.Inst_controller.n8486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i3_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22801\,
            in1 => \N__22849\,
            in2 => \_gnd_net_\,
            in3 => \N__22421\,
            lcout => \syncedInput_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i0_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22325\,
            in1 => \N__22802\,
            in2 => \_gnd_net_\,
            in3 => \N__22622\,
            lcout => \syncedInput_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i5_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29482\,
            in1 => \N__24823\,
            in2 => \_gnd_net_\,
            in3 => \N__31370\,
            lcout => \valueRegister_5_adj_1331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i7_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22477\,
            in1 => \N__29483\,
            in2 => \_gnd_net_\,
            in3 => \N__27199\,
            lcout => \valueRegister_7_adj_1329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27050\,
            in1 => \N__35984\,
            in2 => \_gnd_net_\,
            in3 => \N__26902\,
            lcout => \maskRegister_0_adj_1328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i3_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31163\,
            in1 => \N__32313\,
            in2 => \N__22502\,
            in3 => \N__31955\,
            lcout => \memoryOut_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i7_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__22951\,
            in1 => \N__22751\,
            in2 => \N__26969\,
            in3 => \N__22874\,
            lcout => \syncedInput_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i7_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100101101100"
        )
    port map (
            in0 => \N__35612\,
            in1 => \N__22478\,
            in2 => \N__25106\,
            in3 => \N__23036\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37571\,
            ce => 'H',
            sr => \N__26456\
        );

    \Inst_core.Inst_sampler.i7222_4_lut_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__25054\,
            in1 => \N__27854\,
            in2 => \N__32056\,
            in3 => \N__27806\,
            lcout => \Inst_core.Inst_sampler.n8590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7234_4_lut_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__31655\,
            in1 => \N__24871\,
            in2 => \N__24899\,
            in3 => \N__27506\,
            lcout => \Inst_core.Inst_sampler.n8602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.i1678_3_lut_4_lut_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__22600\,
            in1 => \N__26359\,
            in2 => \N__22466\,
            in3 => \N__23276\,
            lcout => \Inst_core.Inst_sync.n2787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.i5524_1_lut_2_lut_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__26358\,
            in1 => \N__22599\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.n2564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.i1682_3_lut_4_lut_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__23204\,
            in1 => \N__22598\,
            in2 => \N__22442\,
            in3 => \N__26360\,
            lcout => \Inst_core.Inst_sync.n2791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.i1684_3_lut_4_lut_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__26361\,
            in1 => \N__22601\,
            in2 => \N__22646\,
            in3 => \N__22661\,
            lcout => \Inst_core.Inst_sync.n2793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.i1459_3_lut_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__22616\,
            in1 => \N__22597\,
            in2 => \_gnd_net_\,
            in3 => \N__26357\,
            lcout => \Inst_core.Inst_sync.n2566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.output_i1_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22559\,
            in1 => \N__22803\,
            in2 => \_gnd_net_\,
            in3 => \N__22535\,
            lcout => \syncedInput_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i5_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22828\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i6_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31138\,
            in1 => \N__30405\,
            in2 => \N__22523\,
            in3 => \N__31949\,
            lcout => \memoryOut_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i15_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33914\,
            in1 => \N__31140\,
            in2 => \_gnd_net_\,
            in3 => \N__24803\,
            lcout => divider_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i6_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22711\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i16_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31137\,
            in1 => \N__36185\,
            in2 => \_gnd_net_\,
            in3 => \N__24749\,
            lcout => divider_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35997\,
            in1 => \N__31139\,
            in2 => \_gnd_net_\,
            in3 => \N__31567\,
            lcout => divider_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_demux.output_7__11_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23203\,
            lcout => \Inst_core.Inst_sync.demuxedInput_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i2_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23261\,
            lcout => \Inst_core.Inst_sync.demuxedInput_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_demux.output_5__13_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23275\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.demuxedInput_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.n2566_bdd_4_lut_7729_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__22752\,
            in1 => \N__22806\,
            in2 => \N__31435\,
            in3 => \N__23110\,
            lcout => \Inst_core.Inst_sync.n9117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i3_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23228\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.demuxedInput_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i5_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23150\,
            lcout => \Inst_core.Inst_sync.synchronizedInput_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.n2566_bdd_4_lut_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__22805\,
            in1 => \N__22753\,
            in2 => \N__22707\,
            in3 => \N__23161\,
            lcout => \Inst_core.Inst_sync.n9129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i6_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.synchronizedInput_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22681\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23303\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i3_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23227\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i6_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23188\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i5_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23149\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput180_i7_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31459\,
            lcout => \Inst_core.Inst_sync.synchronizedInput180_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVInst_core.Inst_sync.synchronizedInput180_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_2_lut_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__36635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25226\,
            lcout => \Inst_core.n8518\,
            ltout => \Inst_core.n8518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_decoder.i17_4_lut_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__23641\,
            in1 => \N__32503\,
            in2 => \N__23099\,
            in3 => \N__32602\,
            lcout => \Inst_core.Inst_decoder.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i7_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101100101101010"
        )
    port map (
            in0 => \N__23096\,
            in1 => \N__30345\,
            in2 => \N__23078\,
            in3 => \N__23054\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37607\,
            ce => 'H',
            sr => \N__26918\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i7501_2_lut_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25227\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36634\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n8808_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_4_lut_adj_73_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__25241\,
            in1 => \N__36854\,
            in2 => \N__23414\,
            in3 => \N__25183\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i7621_2_lut_3_lut_4_lut_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__25228\,
            in1 => \N__36636\,
            in2 => \N__36873\,
            in3 => \N__25184\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i2_3_lut_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36633\,
            in1 => \N__25182\,
            in2 => \_gnd_net_\,
            in3 => \N__25225\,
            lcout => \Inst_core.n1639\,
            ltout => \Inst_core.n1639_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7669_1_lut_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23405\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.n9054\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i0_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__28136\,
            in1 => \N__23402\,
            in2 => \N__23396\,
            in3 => \N__23381\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7899\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i1_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23378\,
            in1 => \N__23363\,
            in2 => \N__23770\,
            in3 => \N__23351\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7899\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7900\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i2_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23348\,
            in1 => \N__23333\,
            in2 => \N__23751\,
            in3 => \N__23321\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7900\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7901\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i3_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__23318\,
            in1 => \N__23721\,
            in2 => \N__23591\,
            in3 => \N__23576\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7901\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7902\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i4_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__25658\,
            in1 => \N__23569\,
            in2 => \N__23752\,
            in3 => \N__23555\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7902\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7903\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i5_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__23867\,
            in1 => \N__23725\,
            in2 => \N__23551\,
            in3 => \N__23531\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7903\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7904\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i6_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24353\,
            in1 => \N__23528\,
            in2 => \N__23753\,
            in3 => \N__23516\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7904\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7905\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i7_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__23618\,
            in1 => \N__23729\,
            in2 => \N__23513\,
            in3 => \N__23495\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7905\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7906\,
            clk => \N__37598\,
            ce => \N__23669\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i8_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__24017\,
            in1 => \N__23492\,
            in2 => \N__23771\,
            in3 => \N__23480\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8\,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7907\,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i9_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__23837\,
            in1 => \N__23757\,
            in2 => \N__23477\,
            in3 => \N__23462\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7907\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7908\,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i10_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23459\,
            in1 => \N__23447\,
            in2 => \N__23772\,
            in3 => \N__23435\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7908\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7909\,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i11_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__23603\,
            in1 => \N__23761\,
            in2 => \N__23432\,
            in3 => \N__23417\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7909\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7910\,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i12_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__25955\,
            in1 => \N__23822\,
            in2 => \N__23773\,
            in3 => \N__23810\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7910\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7911\,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i13_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__25562\,
            in1 => \N__23765\,
            in2 => \N__23807\,
            in3 => \N__23792\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7911\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7912\,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i14_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23852\,
            in1 => \N__23789\,
            in2 => \N__23774\,
            in3 => \N__23777\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7912\,
            carryout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7913\,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i15_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__23769\,
            in1 => \N__23683\,
            in2 => \N__23939\,
            in3 => \N__23687\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37587\,
            ce => \N__23668\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i25_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23640\,
            in1 => \N__28178\,
            in2 => \_gnd_net_\,
            in3 => \N__35856\,
            lcout => \Inst_core.configRegister_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i14_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29354\,
            in1 => \N__34810\,
            in2 => \N__30119\,
            in3 => \N__35069\,
            lcout => cmd_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i8_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27197\,
            in1 => \N__23614\,
            in2 => \_gnd_net_\,
            in3 => \N__35857\,
            lcout => \configRegister_7_adj_1353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i12_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35854\,
            in1 => \N__34591\,
            in2 => \_gnd_net_\,
            in3 => \N__23602\,
            lcout => \configRegister_11_adj_1349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i13_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26136\,
            in1 => \N__35308\,
            in2 => \_gnd_net_\,
            in3 => \N__23878\,
            lcout => \configRegister_12_adj_1388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i6_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35855\,
            in1 => \N__31374\,
            in2 => \_gnd_net_\,
            in3 => \N__23863\,
            lcout => \configRegister_5_adj_1355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i3_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32749\,
            in1 => \N__34121\,
            in2 => \_gnd_net_\,
            in3 => \N__29678\,
            lcout => \configRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i3_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36104\,
            in1 => \N__26698\,
            in2 => \_gnd_net_\,
            in3 => \N__32392\,
            lcout => \valueRegister_3_adj_1373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i4_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34123\,
            in1 => \N__32719\,
            in2 => \_gnd_net_\,
            in3 => \N__26654\,
            lcout => \configRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i15_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35852\,
            in1 => \N__30114\,
            in2 => \_gnd_net_\,
            in3 => \N__23848\,
            lcout => \configRegister_14_adj_1346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i11_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34122\,
            in1 => \N__25593\,
            in2 => \_gnd_net_\,
            in3 => \N__33076\,
            lcout => \configRegister_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i13_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29310\,
            in1 => \N__35307\,
            in2 => \_gnd_net_\,
            in3 => \N__28372\,
            lcout => \configRegister_12_adj_1308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i10_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23833\,
            in1 => \N__35813\,
            in2 => \_gnd_net_\,
            in3 => \N__26597\,
            lcout => \configRegister_9_adj_1351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i8_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29311\,
            in1 => \N__28507\,
            in2 => \_gnd_net_\,
            in3 => \N__27192\,
            lcout => \configRegister_7_adj_1313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i9_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35853\,
            in1 => \N__24010\,
            in2 => \_gnd_net_\,
            in3 => \N__23999\,
            lcout => \configRegister_8_adj_1352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i18_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29555\,
            in1 => \N__35851\,
            in2 => \_gnd_net_\,
            in3 => \N__28927\,
            lcout => \configRegister_17_adj_1343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i9_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34095\,
            in1 => \N__33130\,
            in2 => \_gnd_net_\,
            in3 => \N__23993\,
            lcout => \configRegister_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i8_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34085\,
            in1 => \N__33163\,
            in2 => \_gnd_net_\,
            in3 => \N__27174\,
            lcout => \configRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23919\,
            in1 => \N__34237\,
            in2 => \_gnd_net_\,
            in3 => \N__26426\,
            lcout => \maskRegister_1_adj_1367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i17_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29554\,
            in1 => \N__31198\,
            in2 => \_gnd_net_\,
            in3 => \N__27237\,
            lcout => divider_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i16_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35850\,
            in1 => \N__33928\,
            in2 => \_gnd_net_\,
            in3 => \N__23932\,
            lcout => \configRegister_15_adj_1345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26441\,
            in1 => \N__35928\,
            in2 => \_gnd_net_\,
            in3 => \N__23918\,
            lcout => \maskRegister_0_adj_1368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i2_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23920\,
            in1 => \N__29677\,
            in2 => \_gnd_net_\,
            in3 => \N__26414\,
            lcout => \maskRegister_2_adj_1366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i11_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29330\,
            in1 => \N__25609\,
            in2 => \_gnd_net_\,
            in3 => \N__28426\,
            lcout => \configRegister_10_adj_1310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i6_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27053\,
            in1 => \N__34420\,
            in2 => \_gnd_net_\,
            in3 => \N__25868\,
            lcout => \maskRegister_6_adj_1322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i13_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29382\,
            in1 => \_gnd_net_\,
            in2 => \N__31199\,
            in3 => \N__24771\,
            lcout => divider_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i5_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27052\,
            in1 => \N__31364\,
            in2 => \_gnd_net_\,
            in3 => \N__25895\,
            lcout => \maskRegister_5_adj_1323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i10_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26585\,
            in1 => \N__26120\,
            in2 => \_gnd_net_\,
            in3 => \N__24073\,
            lcout => \configRegister_9_adj_1391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i24_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35671\,
            in1 => \_gnd_net_\,
            in2 => \N__26135\,
            in3 => \N__33514\,
            lcout => \configRegister_26_adj_1377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i10_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35444\,
            in1 => \N__25608\,
            in2 => \_gnd_net_\,
            in3 => \N__24463\,
            lcout => bwd_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i14_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31192\,
            in2 => \N__30113\,
            in3 => \N__24711\,
            lcout => divider_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i14_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24062\,
            in1 => \N__24034\,
            in2 => \_gnd_net_\,
            in3 => \N__35478\,
            lcout => \Inst_core.Inst_controller.fwd_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i23_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__34960\,
            in1 => \N__29752\,
            in2 => \N__24168\,
            in3 => \N__34789\,
            lcout => cmd_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i10_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__26584\,
            in1 => \N__34961\,
            in2 => \N__25613\,
            in3 => \N__34802\,
            lcout => cmd_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i18_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29541\,
            in1 => \N__26127\,
            in2 => \_gnd_net_\,
            in3 => \N__25801\,
            lcout => \configRegister_17_adj_1383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i26_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__24099\,
            in1 => \N__34962\,
            in2 => \N__34826\,
            in3 => \N__35672\,
            lcout => cmd_33,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i11_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35477\,
            in1 => \N__34592\,
            in2 => \_gnd_net_\,
            in3 => \N__24283\,
            lcout => bwd_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i28_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__24371\,
            in1 => \N__34963\,
            in2 => \N__28176\,
            in3 => \N__34803\,
            lcout => cmd_35,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i21_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24152\,
            in1 => \_gnd_net_\,
            in2 => \N__34119\,
            in3 => \N__24117\,
            lcout => \configRegister_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i4_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29114\,
            in1 => \N__26752\,
            in2 => \_gnd_net_\,
            in3 => \N__35510\,
            lcout => bwd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35509\,
            in1 => \_gnd_net_\,
            in2 => \N__29691\,
            in3 => \N__29932\,
            lcout => bwd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i29_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__34799\,
            in1 => \N__35053\,
            in2 => \N__24395\,
            in3 => \N__24366\,
            lcout => cmd_36,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i9_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35514\,
            in1 => \N__24100\,
            in2 => \_gnd_net_\,
            in3 => \N__24199\,
            lcout => fwd_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i13_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24391\,
            in1 => \N__35512\,
            in2 => \_gnd_net_\,
            in3 => \N__24212\,
            lcout => fwd_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35513\,
            in1 => \N__29540\,
            in2 => \_gnd_net_\,
            in3 => \N__24484\,
            lcout => fwd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i12_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24502\,
            in1 => \N__24367\,
            in2 => \_gnd_net_\,
            in3 => \N__35511\,
            lcout => fwd_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35831\,
            in1 => \N__24346\,
            in2 => \_gnd_net_\,
            in3 => \N__34423\,
            lcout => \configRegister_6_adj_1354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i5_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001011010"
        )
    port map (
            in0 => \N__24335\,
            in1 => \N__24317\,
            in2 => \N__25514\,
            in3 => \N__30332\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37547\,
            ce => 'H',
            sr => \N__24296\
        );

    \Inst_core.Inst_controller.i2_4_lut_adj_60_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__37772\,
            in1 => \N__24284\,
            in2 => \N__24269\,
            in3 => \N__36929\,
            lcout => \Inst_core.Inst_controller.n18_adj_990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i6_4_lut_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24250\,
            in1 => \N__37078\,
            in2 => \N__26486\,
            in3 => \N__37771\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_controller.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i9_4_lut_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__24235\,
            in1 => \N__37051\,
            in2 => \N__24221\,
            in3 => \N__24422\,
            lcout => \Inst_core.Inst_controller.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i3_4_lut_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24211\,
            in1 => \N__36901\,
            in2 => \N__24200\,
            in3 => \N__37724\,
            lcout => \Inst_core.Inst_controller.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i4_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010110101111000"
        )
    port map (
            in0 => \N__30358\,
            in1 => \N__24587\,
            in2 => \N__24560\,
            in3 => \N__28085\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37559\,
            ce => 'H',
            sr => \N__24539\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_adj_71_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24527\,
            in1 => \N__30233\,
            in2 => \N__24521\,
            in3 => \N__24509\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i1_4_lut_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24503\,
            in1 => \N__36211\,
            in2 => \N__24488\,
            in3 => \N__37747\,
            lcout => \Inst_core.Inst_controller.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i4_4_lut_adj_59_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37748\,
            in1 => \N__24464\,
            in2 => \N__35240\,
            in3 => \N__37796\,
            lcout => \Inst_core.Inst_controller.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i8_4_lut_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__34142\,
            in1 => \N__36953\,
            in2 => \N__36215\,
            in3 => \N__27076\,
            lcout => \Inst_core.Inst_controller.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i2_4_lut_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__36952\,
            in1 => \N__27064\,
            in2 => \N__28985\,
            in3 => \N__37795\,
            lcout => \Inst_core.Inst_controller.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.counter_17__I_0_43_i11_2_lut_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24443\,
            in2 => \_gnd_net_\,
            in3 => \N__36928\,
            lcout => \Inst_core.Inst_controller.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register_80_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100010001"
        )
    port map (
            in0 => \N__24416\,
            in1 => \N__24401\,
            in2 => \_gnd_net_\,
            in3 => \N__26362\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27051\,
            in1 => \N__34257\,
            in2 => \_gnd_net_\,
            in3 => \N__27476\,
            lcout => \maskRegister_1_adj_1327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i21_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24686\,
            in1 => \N__31168\,
            in2 => \_gnd_net_\,
            in3 => \N__25027\,
            lcout => divider_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__31166\,
            in1 => \N__24635\,
            in2 => \N__31788\,
            in3 => \N__31953\,
            lcout => \memoryOut_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i4_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29494\,
            in1 => \N__24607\,
            in2 => \_gnd_net_\,
            in3 => \N__29132\,
            lcout => \valueRegister_4_adj_1332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3597_1_lut_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34258\,
            in1 => \_gnd_net_\,
            in2 => \N__29495\,
            in3 => \N__25066\,
            lcout => \valueRegister_1_adj_1335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.sample_i0_i1_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31167\,
            in1 => \N__33608\,
            in2 => \N__24629\,
            in3 => \N__31954\,
            lcout => \memoryOut_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i4_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__25145\,
            in1 => \N__35606\,
            in2 => \N__24614\,
            in3 => \N__28072\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37586\,
            ce => 'H',
            sr => \N__24596\
        );

    \Inst_core.Inst_sampler.i7_4_lut_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__25023\,
            in1 => \N__27850\,
            in2 => \N__29971\,
            in3 => \N__27805\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sampler.n31_adj_995_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i20_4_lut_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24731\,
            in1 => \N__27332\,
            in2 => \N__24590\,
            in3 => \N__24848\,
            lcout => \Inst_core.Inst_sampler.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i5_4_lut_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24895\,
            in1 => \N__27525\,
            in2 => \N__24872\,
            in3 => \N__27701\,
            lcout => \Inst_core.Inst_sampler.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_adj_72_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27383\,
            in1 => \N__24842\,
            in2 => \N__24812\,
            in3 => \N__24833\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7_adj_996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i5_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011111011000"
        )
    port map (
            in0 => \N__35601\,
            in1 => \N__25124\,
            in2 => \N__25511\,
            in3 => \N__24827\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37597\,
            ce => 'H',
            sr => \N__25883\
        );

    \Inst_core.Inst_sampler.i4_4_lut_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24801\,
            in1 => \N__27648\,
            in2 => \N__24778\,
            in3 => \N__27612\,
            lcout => \Inst_core.Inst_sampler.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7236_4_lut_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__24802\,
            in1 => \N__27631\,
            in2 => \N__24785\,
            in3 => \N__31548\,
            lcout => \Inst_core.Inst_sampler.n8604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7230_4_lut_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__24748\,
            in1 => \N__27613\,
            in2 => \N__29975\,
            in3 => \N__30617\,
            lcout => \Inst_core.Inst_sampler.n8598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i8_4_lut_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24747\,
            in1 => \N__27630\,
            in2 => \N__24724\,
            in3 => \N__27592\,
            lcout => \Inst_core.Inst_sampler.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7228_4_lut_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__27299\,
            in1 => \N__27649\,
            in2 => \N__24725\,
            in3 => \N__27699\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sampler.n8596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7300_4_lut_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27215\,
            in1 => \N__27326\,
            in2 => \N__24695\,
            in3 => \N__24692\,
            lcout => \Inst_core.Inst_sampler.n8669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110010101101010"
        )
    port map (
            in0 => \N__25070\,
            in1 => \N__24914\,
            in2 => \N__35611\,
            in3 => \N__33633\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37606\,
            ce => 'H',
            sr => \N__27464\
        );

    \Inst_core.Inst_sampler.i11_4_lut_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__25055\,
            in1 => \N__27876\,
            in2 => \N__27248\,
            in3 => \N__27822\,
            lcout => \Inst_core.Inst_sampler.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7232_4_lut_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__27823\,
            in1 => \N__27362\,
            in2 => \N__25031\,
            in3 => \N__30501\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sampler.n8600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7302_4_lut_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25007\,
            in1 => \N__24998\,
            in2 => \N__24989\,
            in3 => \N__24986\,
            lcout => \Inst_core.Inst_sampler.n8671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i0_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__26390\,
            in1 => \N__24937\,
            in2 => \N__24980\,
            in3 => \N__24956\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24938\,
            in1 => \N__32190\,
            in2 => \_gnd_net_\,
            in3 => \N__26383\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i2_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26384\,
            in1 => \_gnd_net_\,
            in2 => \N__32197\,
            in3 => \N__24912\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i3_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24913\,
            in1 => \N__30816\,
            in2 => \_gnd_net_\,
            in3 => \N__26385\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i4_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26386\,
            in1 => \_gnd_net_\,
            in2 => \N__30823\,
            in3 => \N__31617\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i5_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31618\,
            in1 => \N__25137\,
            in2 => \_gnd_net_\,
            in3 => \N__26387\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i6_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26388\,
            in1 => \_gnd_net_\,
            in2 => \N__25144\,
            in3 => \N__25119\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i7_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25120\,
            in1 => \N__27415\,
            in2 => \_gnd_net_\,
            in3 => \N__26389\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i7564_4_lut_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__25365\,
            in1 => \N__27723\,
            in2 => \N__36657\,
            in3 => \N__25746\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n8844_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.run_83_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36859\,
            in1 => \_gnd_net_\,
            in2 => \N__25091\,
            in3 => \N__32524\,
            lcout => \Inst_core.Inst_trigger.stageRun_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.run_83_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__32440\,
            in1 => \N__36860\,
            in2 => \_gnd_net_\,
            in3 => \N__32555\,
            lcout => \Inst_core.Inst_trigger.stageRun_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.run_83_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__25185\,
            in1 => \_gnd_net_\,
            in2 => \N__36874\,
            in3 => \N__25088\,
            lcout => \Inst_core.stageRun_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i7644_4_lut_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__25366\,
            in1 => \N__25745\,
            in2 => \N__36656\,
            in3 => \N__36858\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n8622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i7667_1_lut_2_lut_3_lut_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__25743\,
            in1 => \N__36625\,
            in2 => \_gnd_net_\,
            in3 => \N__25363\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n9052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i25_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26106\,
            in1 => \N__28199\,
            in2 => \_gnd_net_\,
            in3 => \N__27724\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i890_2_lut_3_lut_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25744\,
            in1 => \N__36626\,
            in2 => \_gnd_net_\,
            in3 => \N__25364\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n1765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i199_2_lut_3_lut_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25204\,
            in1 => \N__26188\,
            in2 => \_gnd_net_\,
            in3 => \N__28879\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n667\,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n667_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i3_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__36663\,
            in1 => \N__25186\,
            in2 => \N__25235\,
            in3 => \N__25232\,
            lcout => \Inst_core.state_1_adj_1134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37609\,
            ce => 'H',
            sr => \N__36865\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i44_2_lut_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26189\,
            in2 => \_gnd_net_\,
            in3 => \N__28880\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i2_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__25154\,
            in1 => \N__25934\,
            in2 => \N__25208\,
            in3 => \N__25205\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37609\,
            ce => 'H',
            sr => \N__36865\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i3_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__28326\,
            in1 => \N__32957\,
            in2 => \N__27911\,
            in3 => \N__36664\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37609\,
            ce => 'H',
            sr => \N__36865\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i1_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__25153\,
            in1 => \N__25196\,
            in2 => \N__25190\,
            in3 => \N__25935\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37609\,
            ce => 'H',
            sr => \N__36865\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i1_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__25932\,
            in1 => \N__25399\,
            in2 => \_gnd_net_\,
            in3 => \N__28358\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37609\,
            ce => 'H',
            sr => \N__36865\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i2_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__25841\,
            in1 => \N__25933\,
            in2 => \N__25403\,
            in3 => \N__25831\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37609\,
            ce => 'H',
            sr => \N__36865\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25739\,
            in2 => \_gnd_net_\,
            in3 => \N__25361\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i1_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__25937\,
            in1 => \N__36646\,
            in2 => \N__25391\,
            in3 => \N__25375\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n760\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \N__36864\
        );

    \Inst_core.Inst_sampler.i1_2_lut_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36645\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32433\,
            lcout => OPEN,
            ltout => \Inst_core.n8515_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i1_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__25939\,
            in1 => \N__25384\,
            in2 => \N__25388\,
            in3 => \N__33268\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \N__36864\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i2_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__25385\,
            in1 => \N__25936\,
            in2 => \N__28573\,
            in3 => \N__28589\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \N__36864\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i2_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__25938\,
            in1 => \N__25376\,
            in2 => \N__25775\,
            in3 => \N__25787\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \N__36864\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i3_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001100"
        )
    port map (
            in0 => \N__33269\,
            in1 => \N__32434\,
            in2 => \N__36662\,
            in3 => \N__32474\,
            lcout => \Inst_core.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \N__36864\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i3_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110110000"
        )
    port map (
            in0 => \N__25362\,
            in1 => \N__36647\,
            in2 => \N__25748\,
            in3 => \N__25757\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \N__36864\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register_80_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100010001"
        )
    port map (
            in0 => \N__32675\,
            in1 => \N__27926\,
            in2 => \_gnd_net_\,
            in3 => \N__26382\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i6_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29252\,
            in1 => \N__28549\,
            in2 => \_gnd_net_\,
            in3 => \N__31383\,
            lcout => \configRegister_5_adj_1315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i10_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25599\,
            in1 => \N__31031\,
            in2 => \_gnd_net_\,
            in3 => \N__27294\,
            lcout => divider_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i4_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29251\,
            in1 => \N__28234\,
            in2 => \_gnd_net_\,
            in3 => \N__26725\,
            lcout => \configRegister_3_adj_1317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i14_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35858\,
            in1 => \N__29355\,
            in2 => \_gnd_net_\,
            in3 => \N__25558\,
            lcout => \configRegister_13_adj_1347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i15_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26137\,
            in1 => \N__30115\,
            in2 => \_gnd_net_\,
            in3 => \N__25543\,
            lcout => \configRegister_14_adj_1386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i7_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34433\,
            in1 => \N__29253\,
            in2 => \_gnd_net_\,
            in3 => \N__28531\,
            lcout => \configRegister_6_adj_1314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i3_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29250\,
            in1 => \N__28255\,
            in2 => \_gnd_net_\,
            in3 => \N__29675\,
            lcout => \configRegister_2_adj_1318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i5_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001011010"
        )
    port map (
            in0 => \N__26177\,
            in1 => \N__25532\,
            in2 => \N__25507\,
            in3 => \N__33551\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37576\,
            ce => 'H',
            sr => \N__25625\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_2_lut_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26612\,
            in2 => \_gnd_net_\,
            in3 => \N__28956\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i44_4_lut_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100000000"
        )
    port map (
            in0 => \N__25673\,
            in1 => \N__28910\,
            in2 => \N__25856\,
            in3 => \N__25853\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n100\,
            ltout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i166_2_lut_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__25832\,
            in1 => \_gnd_net_\,
            in2 => \N__25817\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_74_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25970\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i44_4_lut_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001100"
        )
    port map (
            in0 => \N__28911\,
            in1 => \N__25814\,
            in2 => \N__25808\,
            in3 => \N__25805\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n100\,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i232_2_lut_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25778\,
            in3 => \N__25774\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n770\,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n770_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_4_lut_adj_75_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__25747\,
            in1 => \N__36808\,
            in2 => \N__25709\,
            in3 => \N__25706\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4076\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i18_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29318\,
            in1 => \N__29548\,
            in2 => \_gnd_net_\,
            in3 => \N__25672\,
            lcout => \configRegister_17_adj_1303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i5_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29122\,
            in1 => \N__35835\,
            in2 => \_gnd_net_\,
            in3 => \N__25651\,
            lcout => \configRegister_4_adj_1356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3605_1_lut_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25640\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i10_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34096\,
            in1 => \N__33109\,
            in2 => \_gnd_net_\,
            in3 => \N__26595\,
            lcout => \configRegister_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i10_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26594\,
            in1 => \N__29320\,
            in2 => \_gnd_net_\,
            in3 => \N__28462\,
            lcout => \configRegister_9_adj_1311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i13_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35289\,
            in1 => \N__35834\,
            in2 => \_gnd_net_\,
            in3 => \N__25951\,
            lcout => \configRegister_12_adj_1348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i5_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29319\,
            in1 => \N__28213\,
            in2 => \_gnd_net_\,
            in3 => \N__29123\,
            lcout => \configRegister_4_adj_1316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i15_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34097\,
            in1 => \N__30100\,
            in2 => \_gnd_net_\,
            in3 => \N__33814\,
            lcout => \configRegister_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.levelReg_927__i1_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__28955\,
            in1 => \_gnd_net_\,
            in2 => \N__33368\,
            in3 => \N__28909\,
            lcout => \Inst_core.Inst_trigger.levelReg_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37549\,
            ce => 'H',
            sr => \N__25940\
        );

    \Inst_core.Inst_trigger.levelReg_927__i0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33364\,
            in2 => \_gnd_net_\,
            in3 => \N__28954\,
            lcout => \Inst_core.Inst_trigger.levelReg_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37549\,
            ce => 'H',
            sr => \N__25940\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3598_1_lut_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25894\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3599_1_lut_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25867\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3600_1_lut_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26471\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3486_1_lut_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26437\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3601_1_lut_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26425\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4760\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3602_1_lut_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26413\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n4761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register_80_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100010001"
        )
    port map (
            in0 => \N__32123\,
            in1 => \N__26402\,
            in2 => \_gnd_net_\,
            in3 => \N__26381\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i5_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31332\,
            in1 => \N__36103\,
            in2 => \_gnd_net_\,
            in3 => \N__26173\,
            lcout => \valueRegister_5_adj_1371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30205\,
            in1 => \N__36175\,
            in2 => \_gnd_net_\,
            in3 => \N__35466\,
            lcout => fwd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i14_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29394\,
            in1 => \N__26144\,
            in2 => \_gnd_net_\,
            in3 => \N__26155\,
            lcout => \configRegister_13_adj_1387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i17_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26143\,
            in1 => \N__36177\,
            in2 => \_gnd_net_\,
            in3 => \N__25969\,
            lcout => \configRegister_16_adj_1384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i17_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36176\,
            in1 => \N__29325\,
            in2 => \_gnd_net_\,
            in3 => \N__26611\,
            lcout => \configRegister_16_adj_1304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i9_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35465\,
            in1 => \N__26587\,
            in2 => \_gnd_net_\,
            in3 => \N__26887\,
            lcout => bwd_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i13_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__35270\,
            in1 => \N__34821\,
            in2 => \N__29399\,
            in3 => \N__35055\,
            lcout => cmd_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i20_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__35054\,
            in1 => \N__26540\,
            in2 => \N__34842\,
            in3 => \N__29988\,
            lcout => cmd_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i6_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35516\,
            in1 => \N__34428\,
            in2 => \_gnd_net_\,
            in3 => \N__26801\,
            lcout => bwd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26729\,
            in1 => \N__29475\,
            in2 => \_gnd_net_\,
            in3 => \N__31594\,
            lcout => \valueRegister_3_adj_1333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27049\,
            in1 => \N__26728\,
            in2 => \_gnd_net_\,
            in3 => \N__27436\,
            lcout => \maskRegister_3_adj_1325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26727\,
            in1 => \N__34521\,
            in2 => \_gnd_net_\,
            in3 => \N__26842\,
            lcout => \valueRegister_3_adj_1293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35515\,
            in1 => \N__26726\,
            in2 => \_gnd_net_\,
            in3 => \N__26765\,
            lcout => bwd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i3_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35517\,
            in1 => \N__29989\,
            in2 => \_gnd_net_\,
            in3 => \N__26485\,
            lcout => fwd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i6_4_lut_adj_58_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__26888\,
            in1 => \N__37664\,
            in2 => \N__28832\,
            in3 => \N__36902\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_controller.n22_adj_988_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i14_4_lut_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26873\,
            in1 => \N__26771\,
            in2 => \N__26867\,
            in3 => \N__26738\,
            lcout => \Inst_core.Inst_controller.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i3_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__26864\,
            in1 => \N__26843\,
            in2 => \N__30346\,
            in3 => \N__32351\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37561\,
            ce => 'H',
            sr => \N__26813\
        );

    \Inst_core.Inst_controller.i7_4_lut_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__26800\,
            in1 => \N__37024\,
            in2 => \N__26789\,
            in3 => \N__36988\,
            lcout => \Inst_core.Inst_controller.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i5_4_lut_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37052\,
            in1 => \N__26764\,
            in2 => \N__26753\,
            in3 => \N__37079\,
            lcout => \Inst_core.Inst_controller.n21_adj_989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i2_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31112\,
            in1 => \N__29713\,
            in2 => \_gnd_net_\,
            in3 => \N__27315\,
            lcout => divider_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i18_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30035\,
            in1 => \N__31114\,
            in2 => \_gnd_net_\,
            in3 => \N__30579\,
            lcout => divider_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31113\,
            in1 => \N__26731\,
            in2 => \_gnd_net_\,
            in3 => \N__31683\,
            lcout => divider_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29711\,
            in1 => \N__27042\,
            in2 => \_gnd_net_\,
            in3 => \N__27449\,
            lcout => \maskRegister_2_adj_1326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i7_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35518\,
            in1 => \N__27207\,
            in2 => \_gnd_net_\,
            in3 => \N__27077\,
            lcout => bwd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29712\,
            in1 => \N__29490\,
            in2 => \_gnd_net_\,
            in3 => \N__30838\,
            lcout => \valueRegister_2_adj_1334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i10_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35519\,
            in1 => \N__35680\,
            in2 => \_gnd_net_\,
            in3 => \N__27065\,
            lcout => fwd_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i4_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27043\,
            in1 => \N__29129\,
            in2 => \_gnd_net_\,
            in3 => \N__26981\,
            lcout => \maskRegister_4_adj_1324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.result_i7_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__26962\,
            in1 => \N__31472\,
            in2 => \_gnd_net_\,
            in3 => \N__31436\,
            lcout => \Inst_core.Inst_sync.filteredInput_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37588\,
            ce => 'H',
            sr => \N__26948\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3593_1_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26936\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i7670_1_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28769\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n9055\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3484_1_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26903\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3594_1_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27475\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3595_1_lut_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27448\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3596_1_lut_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27437\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n4755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i6_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010111001010"
        )
    port map (
            in0 => \N__30452\,
            in1 => \N__27422\,
            in2 => \N__35600\,
            in3 => \N__27404\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37599\,
            ce => 'H',
            sr => \N__27377\
        );

    \Inst_core.Inst_sampler.i6_4_lut_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__30699\,
            in1 => \N__27316\,
            in2 => \N__27361\,
            in3 => \N__27552\,
            lcout => \Inst_core.Inst_sampler.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7224_4_lut_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__27274\,
            in1 => \N__27553\,
            in2 => \N__32108\,
            in3 => \N__27526\,
            lcout => \Inst_core.Inst_sampler.n8592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7238_4_lut_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__30583\,
            in1 => \N__30555\,
            in2 => \N__27887\,
            in3 => \N__27317\,
            lcout => \Inst_core.Inst_sampler.n8606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i9_4_lut_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__27295\,
            in1 => \N__27502\,
            in2 => \N__27275\,
            in3 => \N__27676\,
            lcout => \Inst_core.Inst_sampler.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7220_4_lut_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__27677\,
            in1 => \N__27247\,
            in2 => \N__27596\,
            in3 => \N__30785\,
            lcout => \Inst_core.Inst_sampler.n8588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.counter_926__i0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31497\,
            in2 => \_gnd_net_\,
            in3 => \N__27566\,
            lcout => \Inst_core.Inst_sampler.counter_0\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \Inst_core.Inst_sampler.n7948\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30557\,
            in2 => \_gnd_net_\,
            in3 => \N__27563\,
            lcout => \Inst_core.Inst_sampler.counter_1\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7948\,
            carryout => \Inst_core.Inst_sampler.n7949\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30703\,
            in2 => \_gnd_net_\,
            in3 => \N__27560\,
            lcout => \Inst_core.Inst_sampler.counter_2\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7949\,
            carryout => \Inst_core.Inst_sampler.n7950\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30503\,
            in2 => \_gnd_net_\,
            in3 => \N__27557\,
            lcout => \Inst_core.Inst_sampler.counter_3\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7950\,
            carryout => \Inst_core.Inst_sampler.n7951\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i4_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27554\,
            in2 => \_gnd_net_\,
            in3 => \N__27536\,
            lcout => \Inst_core.Inst_sampler.counter_4\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7951\,
            carryout => \Inst_core.Inst_sampler.n7952\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i5_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32019\,
            in2 => \_gnd_net_\,
            in3 => \N__27533\,
            lcout => \Inst_core.Inst_sampler.counter_5\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7952\,
            carryout => \Inst_core.Inst_sampler.n7953\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i6_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31654\,
            in2 => \_gnd_net_\,
            in3 => \N__27530\,
            lcout => \Inst_core.Inst_sampler.counter_6\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7953\,
            carryout => \Inst_core.Inst_sampler.n7954\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i7_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27527\,
            in2 => \_gnd_net_\,
            in3 => \N__27509\,
            lcout => \Inst_core.Inst_sampler.counter_7\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7954\,
            carryout => \Inst_core.Inst_sampler.n7955\,
            clk => \N__37608\,
            ce => 'H',
            sr => \N__27756\
        );

    \Inst_core.Inst_sampler.counter_926__i8_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27501\,
            in2 => \_gnd_net_\,
            in3 => \N__27479\,
            lcout => \Inst_core.Inst_sampler.counter_8\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \Inst_core.Inst_sampler.n7956\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i9_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27700\,
            in2 => \_gnd_net_\,
            in3 => \N__27680\,
            lcout => \Inst_core.Inst_sampler.counter_9\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7956\,
            carryout => \Inst_core.Inst_sampler.n7957\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i10_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27675\,
            in2 => \_gnd_net_\,
            in3 => \N__27659\,
            lcout => \Inst_core.Inst_sampler.counter_10\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7957\,
            carryout => \Inst_core.Inst_sampler.n7958\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i11_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30721\,
            in2 => \_gnd_net_\,
            in3 => \N__27656\,
            lcout => \Inst_core.Inst_sampler.counter_11\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7958\,
            carryout => \Inst_core.Inst_sampler.n7959\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i12_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31549\,
            in2 => \_gnd_net_\,
            in3 => \N__27653\,
            lcout => \Inst_core.Inst_sampler.counter_12\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7959\,
            carryout => \Inst_core.Inst_sampler.n7960\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i13_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27650\,
            in2 => \_gnd_net_\,
            in3 => \N__27635\,
            lcout => \Inst_core.Inst_sampler.counter_13\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7960\,
            carryout => \Inst_core.Inst_sampler.n7961\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i14_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27632\,
            in2 => \_gnd_net_\,
            in3 => \N__27617\,
            lcout => \Inst_core.Inst_sampler.counter_14\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7961\,
            carryout => \Inst_core.Inst_sampler.n7962\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i15_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27614\,
            in2 => \_gnd_net_\,
            in3 => \N__27599\,
            lcout => \Inst_core.Inst_sampler.counter_15\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7962\,
            carryout => \Inst_core.Inst_sampler.n7963\,
            clk => \N__37615\,
            ce => 'H',
            sr => \N__27763\
        );

    \Inst_core.Inst_sampler.counter_926__i16_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27591\,
            in2 => \_gnd_net_\,
            in3 => \N__27569\,
            lcout => \Inst_core.Inst_sampler.counter_16\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \Inst_core.Inst_sampler.n7964\,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_sampler.counter_926__i17_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27880\,
            in2 => \_gnd_net_\,
            in3 => \N__27860\,
            lcout => \Inst_core.Inst_sampler.counter_17\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7964\,
            carryout => \Inst_core.Inst_sampler.n7965\,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_sampler.counter_926__i18_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30609\,
            in2 => \_gnd_net_\,
            in3 => \N__27857\,
            lcout => \Inst_core.Inst_sampler.counter_18\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7965\,
            carryout => \Inst_core.Inst_sampler.n7966\,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_sampler.counter_926__i19_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27849\,
            in2 => \_gnd_net_\,
            in3 => \N__27827\,
            lcout => \Inst_core.Inst_sampler.counter_19\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7966\,
            carryout => \Inst_core.Inst_sampler.n7967\,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_sampler.counter_926__i20_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27824\,
            in2 => \_gnd_net_\,
            in3 => \N__27809\,
            lcout => \Inst_core.Inst_sampler.counter_20\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7967\,
            carryout => \Inst_core.Inst_sampler.n7968\,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_sampler.counter_926__i21_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27798\,
            in2 => \_gnd_net_\,
            in3 => \N__27776\,
            lcout => \Inst_core.Inst_sampler.counter_21\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7968\,
            carryout => \Inst_core.Inst_sampler.n7969\,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_sampler.counter_926__i22_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32080\,
            in2 => \_gnd_net_\,
            in3 => \N__27773\,
            lcout => \Inst_core.Inst_sampler.counter_22\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_sampler.n7969\,
            carryout => \Inst_core.Inst_sampler.n7970\,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_sampler.counter_926__i23_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30745\,
            in2 => \_gnd_net_\,
            in3 => \N__27770\,
            lcout => \Inst_core.Inst_sampler.counter_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37622\,
            ce => 'H',
            sr => \N__27767\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.match_84_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27728\,
            lcout => \Inst_core.Inst_trigger.stageMatch_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37624\,
            ce => \N__32632\,
            sr => \N__27710\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.run_83_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__32631\,
            in1 => \N__32489\,
            in2 => \N__31862\,
            in3 => \N__28351\,
            lcout => \Inst_core.stageRun_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i25_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28191\,
            in1 => \_gnd_net_\,
            in2 => \N__29324\,
            in3 => \N__31857\,
            lcout => \Inst_core.configRegister_27_adj_1196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i25_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28190\,
            in1 => \N__34105\,
            in2 => \_gnd_net_\,
            in3 => \N__32661\,
            lcout => \Inst_core.Inst_trigger.configRegister_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i1_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29294\,
            in1 => \N__35998\,
            in2 => \_gnd_net_\,
            in3 => \N__28309\,
            lcout => \configRegister_0_adj_1320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i1_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35999\,
            in1 => \N__35833\,
            in2 => \_gnd_net_\,
            in3 => \N__28132\,
            lcout => \configRegister_0_adj_1360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i2_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29295\,
            in1 => \N__34268\,
            in2 => \_gnd_net_\,
            in3 => \N__28270\,
            lcout => \configRegister_1_adj_1319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i4_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011111011000"
        )
    port map (
            in0 => \N__33556\,
            in1 => \N__28121\,
            in2 => \N__28097\,
            in3 => \N__28865\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37611\,
            ce => 'H',
            sr => \N__27986\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_adj_77_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27968\,
            in1 => \N__27956\,
            in2 => \N__27947\,
            in3 => \N__27932\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i5511_2_lut_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36563\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n6675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_4_lut_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__36844\,
            in1 => \N__28339\,
            in2 => \N__27914\,
            in3 => \N__27910\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i12_4_lut_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28789\,
            in1 => \N__28451\,
            in2 => \N__28679\,
            in3 => \N__28394\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i7651_2_lut_4_lut_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__36564\,
            in1 => \N__28338\,
            in2 => \N__36867\,
            in3 => \N__32950\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n8626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i7561_2_lut_3_lut_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__32949\,
            in1 => \N__36565\,
            in2 => \_gnd_net_\,
            in3 => \N__28340\,
            lcout => \Inst_core.n8837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i834_2_lut_3_lut_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36562\,
            in1 => \N__28337\,
            in2 => \_gnd_net_\,
            in3 => \N__32947\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n1662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__28310\,
            in1 => \N__28295\,
            in2 => \N__33014\,
            in3 => \N__28280\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0\,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7884\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i1_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__28277\,
            in1 => \N__28710\,
            in2 => \N__32981\,
            in3 => \N__28259\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7884\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7885\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__28256\,
            in1 => \N__32912\,
            in2 => \N__28743\,
            in3 => \N__28241\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7885\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7886\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i3_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__28238\,
            in1 => \N__28714\,
            in2 => \N__32858\,
            in3 => \N__28223\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7886\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7887\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i4_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__28220\,
            in1 => \N__32995\,
            in2 => \N__28744\,
            in3 => \N__28202\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7887\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7888\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i5_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__28553\,
            in1 => \N__28718\,
            in2 => \N__32831\,
            in3 => \N__28538\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7888\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7889\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i6_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__28535\,
            in1 => \N__32240\,
            in2 => \N__28745\,
            in3 => \N__28520\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7889\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7890\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i7_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__28517\,
            in1 => \N__28722\,
            in2 => \N__32897\,
            in3 => \N__28496\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7890\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7891\,
            clk => \N__37602\,
            ce => \N__28657\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i8_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__28493\,
            in1 => \N__28749\,
            in2 => \N__32813\,
            in3 => \N__28472\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8\,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7892\,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i9_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__28469\,
            in1 => \N__28450\,
            in2 => \N__28766\,
            in3 => \N__28436\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7892\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7893\,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i10_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__28433\,
            in1 => \N__28753\,
            in2 => \N__32879\,
            in3 => \N__28415\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7893\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7894\,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i11_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__28412\,
            in1 => \N__28393\,
            in2 => \N__28767\,
            in3 => \N__28379\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7894\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7895\,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i12_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__28376\,
            in1 => \N__28757\,
            in2 => \N__32930\,
            in3 => \N__28361\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7895\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7896\,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i13_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__28811\,
            in1 => \N__32843\,
            in2 => \N__28768\,
            in3 => \N__28793\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7896\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7897\,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i14_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__29147\,
            in1 => \N__28761\,
            in2 => \N__28790\,
            in3 => \N__28772\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7897\,
            carryout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n7898\,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i15_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__28762\,
            in1 => \N__28675\,
            in2 => \N__28850\,
            in3 => \N__28682\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37591\,
            ce => \N__28661\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i2_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__28646\,
            in1 => \N__33552\,
            in2 => \N__29573\,
            in3 => \N__30928\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37578\,
            ce => 'H',
            sr => \N__28622\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i11_4_lut_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33859\,
            in1 => \N__32737\,
            in2 => \N__33151\,
            in3 => \N__33061\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i12_4_lut_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33799\,
            in1 => \N__33097\,
            in2 => \N__33709\,
            in3 => \N__33028\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_2_lut_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__35084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28963\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i44_4_lut_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100000000"
        )
    port map (
            in0 => \N__29414\,
            in1 => \N__28913\,
            in2 => \N__28607\,
            in3 => \N__28604\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n100\,
            ltout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i133_2_lut_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28577\,
            in3 => \N__28574\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.LessThan_42_i4_4_lut_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28964\,
            in1 => \N__28928\,
            in2 => \N__36125\,
            in3 => \N__28912\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i4_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29130\,
            in1 => \N__28861\,
            in2 => \_gnd_net_\,
            in3 => \N__36092\,
            lcout => \valueRegister_4_adj_1372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i6_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34100\,
            in1 => \N__33202\,
            in2 => \_gnd_net_\,
            in3 => \N__31322\,
            lcout => \configRegister_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i12_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35310\,
            in1 => \N__31091\,
            in2 => \_gnd_net_\,
            in3 => \N__31524\,
            lcout => divider_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34099\,
            in1 => \N__35957\,
            in2 => \_gnd_net_\,
            in3 => \N__32788\,
            lcout => \configRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i16_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29292\,
            in1 => \N__33936\,
            in2 => \_gnd_net_\,
            in3 => \N__28843\,
            lcout => \configRegister_15_adj_1305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i7_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34101\,
            in1 => \N__33184\,
            in2 => \_gnd_net_\,
            in3 => \N__34421\,
            lcout => \configRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i15_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35432\,
            in1 => \N__33935\,
            in2 => \_gnd_net_\,
            in3 => \N__28825\,
            lcout => bwd_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i24_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29293\,
            in1 => \N__30296\,
            in2 => \_gnd_net_\,
            in3 => \N__35676\,
            lcout => \configRegister_26_adj_1297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i18_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29528\,
            in1 => \N__34104\,
            in2 => \_gnd_net_\,
            in3 => \N__29413\,
            lcout => \configRegister_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i13_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29395\,
            in1 => \N__35433\,
            in2 => \_gnd_net_\,
            in3 => \N__29914\,
            lcout => bwd_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34528\,
            in1 => \N__29692\,
            in2 => \_gnd_net_\,
            in3 => \N__29824\,
            lcout => \valueRegister_2_adj_1294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i12_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34102\,
            in1 => \N__34569\,
            in2 => \_gnd_net_\,
            in3 => \N__33040\,
            lcout => \configRegister_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i15_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29143\,
            in1 => \N__29291\,
            in2 => \_gnd_net_\,
            in3 => \N__30085\,
            lcout => \configRegister_14_adj_1306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i5_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34103\,
            in1 => \N__33220\,
            in2 => \_gnd_net_\,
            in3 => \N__29131\,
            lcout => \configRegister_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i6_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34430\,
            in1 => \N__31092\,
            in2 => \_gnd_net_\,
            in3 => \N__30522\,
            lcout => divider_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36099\,
            in1 => \N__34259\,
            in2 => \_gnd_net_\,
            in3 => \N__33664\,
            lcout => \valueRegister_1_adj_1375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i14_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35506\,
            in1 => \N__30069\,
            in2 => \_gnd_net_\,
            in3 => \N__29848\,
            lcout => \Inst_core.Inst_controller.bwd_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i7_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35507\,
            in1 => \N__29764\,
            in2 => \_gnd_net_\,
            in3 => \N__28978\,
            lcout => fwd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i1_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34262\,
            in1 => \N__31090\,
            in2 => \_gnd_net_\,
            in3 => \N__30636\,
            lcout => divider_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i6_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__34431\,
            in1 => \N__34825\,
            in2 => \N__31324\,
            in3 => \N__35052\,
            lcout => cmd_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i3592_1_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29780\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n4751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i23_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31089\,
            in1 => \N__29765\,
            in2 => \_gnd_net_\,
            in3 => \N__30666\,
            lcout => divider_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i2_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36090\,
            in1 => \N__29671\,
            in2 => \_gnd_net_\,
            in3 => \N__29566\,
            lcout => \valueRegister_2_adj_1374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i19_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__35048\,
            in1 => \N__30001\,
            in2 => \N__30034\,
            in3 => \N__34846\,
            lcout => cmd_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i18_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__34843\,
            in1 => \N__29513\,
            in2 => \N__30033\,
            in3 => \N__35049\,
            lcout => cmd_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i17_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__35047\,
            in1 => \N__36146\,
            in2 => \N__29527\,
            in3 => \N__34845\,
            lcout => cmd_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29489\,
            in1 => \N__35989\,
            in2 => \_gnd_net_\,
            in3 => \N__32209\,
            lcout => \valueRegister_0_adj_1336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i15_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__35046\,
            in1 => \N__30068\,
            in2 => \N__33941\,
            in3 => \N__34844\,
            lcout => cmd_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.fwd_i0_i2_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30023\,
            in1 => \N__35508\,
            in2 => \_gnd_net_\,
            in3 => \N__30187\,
            lcout => fwd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i19_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31093\,
            in1 => \_gnd_net_\,
            in2 => \N__30002\,
            in3 => \N__29958\,
            lcout => divider_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i1_4_lut_adj_62_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37723\,
            in1 => \N__29936\,
            in2 => \N__29918\,
            in3 => \N__37099\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_controller.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i13_4_lut_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29900\,
            in1 => \N__29888\,
            in2 => \N__29879\,
            in3 => \N__29834\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_controller.n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i1_3_lut_4_lut_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__36274\,
            in1 => \N__29876\,
            in2 => \N__29864\,
            in3 => \N__36256\,
            lcout => \Inst_core.Inst_controller.nstate_1_N_827_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i5529_2_lut_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36255\,
            in2 => \_gnd_net_\,
            in3 => \N__36273\,
            lcout => \Inst_core.Inst_controller.n6693\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i3_4_lut_adj_61_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__29849\,
            in1 => \N__37696\,
            in2 => \N__35873\,
            in3 => \N__36235\,
            lcout => \Inst_core.Inst_controller.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001011010"
        )
    port map (
            in0 => \N__29828\,
            in1 => \N__29813\,
            in2 => \N__30941\,
            in3 => \N__30344\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37590\,
            ce => 'H',
            sr => \N__30482\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i6_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011011000110"
        )
    port map (
            in0 => \N__30442\,
            in1 => \N__34301\,
            in2 => \N__30347\,
            in3 => \N__30254\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37601\,
            ce => 'H',
            sr => \N__30221\
        );

    \Inst_core.Inst_controller.i4_4_lut_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__30209\,
            in1 => \N__37098\,
            in2 => \N__30191\,
            in3 => \N__36234\,
            lcout => \Inst_core.Inst_controller.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i102_2_lut_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36447\,
            in2 => \_gnd_net_\,
            in3 => \N__36317\,
            lcout => debugleds_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_decoder.i1_2_lut_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__36448\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36871\,
            lcout => OPEN,
            ltout => \Inst_core.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i7628_4_lut_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__36512\,
            in1 => \N__30144\,
            in2 => \N__30125\,
            in3 => \N__36674\,
            lcout => \Inst_core.Inst_controller.n3907\,
            ltout => \Inst_core.Inst_controller.n3907_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i7641_4_lut_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110000"
        )
    port map (
            in0 => \N__36318\,
            in1 => \N__35184\,
            in2 => \N__30122\,
            in3 => \N__36281\,
            lcout => \Inst_core.Inst_controller.n4691\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i7666_3_lut_4_lut_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__33267\,
            in1 => \N__32450\,
            in2 => \N__36553\,
            in3 => \N__36872\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7668_1_lut_2_lut_3_lut_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__32449\,
            in1 => \N__36508\,
            in2 => \_gnd_net_\,
            in3 => \N__33266\,
            lcout => \Inst_core.n9053\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i2_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011011000110"
        )
    port map (
            in0 => \N__30940\,
            in1 => \N__30845\,
            in2 => \N__35578\,
            in3 => \N__30827\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37610\,
            ce => 'H',
            sr => \N__30803\
        );

    \Inst_core.Inst_sampler.i12_4_lut_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__30784\,
            in1 => \N__30727\,
            in2 => \N__30671\,
            in3 => \N__30749\,
            lcout => \Inst_core.Inst_sampler.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7250_4_lut_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__31505\,
            in1 => \N__30638\,
            in2 => \N__30731\,
            in3 => \N__31528\,
            lcout => \Inst_core.Inst_sampler.n8618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.counter_22__I_0_i3_2_lut_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30707\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sampler.n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7288_4_lut_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111110"
        )
    port map (
            in0 => \N__30683\,
            in1 => \N__30524\,
            in2 => \N__30674\,
            in3 => \N__32027\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sampler.n8656_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7304_4_lut_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__30670\,
            in1 => \N__30650\,
            in2 => \N__30641\,
            in3 => \N__32081\,
            lcout => \Inst_core.Inst_sampler.n8673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i3_4_lut_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__30637\,
            in1 => \N__30616\,
            in2 => \N__30590\,
            in3 => \N__30556\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_sampler.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i19_4_lut_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30536\,
            in1 => \N__31631\,
            in2 => \N__30527\,
            in3 => \N__31478\,
            lcout => \Inst_core.Inst_sampler.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i2_4_lut_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__30523\,
            in1 => \N__30502\,
            in2 => \N__31688\,
            in3 => \N__31650\,
            lcout => \Inst_core.Inst_sampler.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__31625\,
            in1 => \N__31604\,
            in2 => \N__35610\,
            in3 => \N__32352\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37617\,
            ce => 'H',
            sr => \N__31583\
        );

    \Inst_core.Inst_sampler.i1_4_lut_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__31568\,
            in1 => \N__31553\,
            in2 => \N__31529\,
            in3 => \N__31498\,
            lcout => \Inst_core.Inst_sampler.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.Inst_filter.input360_i7_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31428\,
            lcout => \Inst_core.Inst_sync.Inst_filter.input360_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sync.synchronizedInput_i7_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Inst_core.Inst_sync.synchronizedInput_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.divider_i0_i5_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31323\,
            in1 => \N__31103\,
            in2 => \_gnd_net_\,
            in3 => \N__32101\,
            lcout => divider_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i21_4_lut_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31997\,
            in1 => \N__31232\,
            in2 => \N__31223\,
            in3 => \N__31211\,
            lcout => \Inst_core.Inst_sampler.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.ready_40_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31102\,
            in2 => \_gnd_net_\,
            in3 => \N__31896\,
            lcout => \sampleReady\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7611_4_lut_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__31895\,
            in1 => \N__30974\,
            in2 => \N__30962\,
            in3 => \N__30950\,
            lcout => \Inst_core.Inst_sampler.n8687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i0_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110010101101010"
        )
    port map (
            in0 => \N__32213\,
            in1 => \N__32198\,
            in2 => \N__35605\,
            in3 => \N__31800\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37627\,
            ce => 'H',
            sr => \N__32177\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32162\,
            in1 => \N__32150\,
            in2 => \N__32141\,
            in3 => \N__32129\,
            lcout => \Inst_core.Inst_trigger.stages_2__Inst_stage.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i10_4_lut_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32097\,
            in1 => \N__32076\,
            in2 => \N__32057\,
            in3 => \N__32026\,
            lcout => \Inst_core.Inst_sampler.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i7609_3_lut_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__31991\,
            in1 => \N__31979\,
            in2 => \_gnd_net_\,
            in3 => \N__31970\,
            lcout => \ready50_N_581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.match_84_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31861\,
            lcout => \Inst_core.Inst_trigger.stageMatch_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37628\,
            ce => \N__32620\,
            sr => \N__31844\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.match_84_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32662\,
            lcout => \Inst_core.Inst_trigger.stageMatch_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37626\,
            ce => \N__32639\,
            sr => \N__31832\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i0_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011010011010"
        )
    port map (
            in0 => \N__36020\,
            in1 => \N__33559\,
            in2 => \N__31804\,
            in3 => \N__31715\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37620\,
            ce => 'H',
            sr => \N__32705\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33443\,
            in1 => \N__32693\,
            in2 => \N__32264\,
            in3 => \N__32681\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7_adj_1000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_76_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__33259\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36612\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n8521_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.i18_4_lut_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__32663\,
            in1 => \N__32542\,
            in2 => \N__32642\,
            in3 => \N__32621\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.i3_4_lut_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32543\,
            in1 => \N__32528\,
            in2 => \N__32510\,
            in3 => \N__32488\,
            lcout => \Inst_core.nstate_1_N_831_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i7508_2_lut_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36611\,
            in2 => \_gnd_net_\,
            in3 => \N__33260\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n8753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_4_lut_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__32439\,
            in1 => \N__36866\,
            in2 => \N__32477\,
            in3 => \N__32473\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n4044\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_sampler.i1_2_lut_3_lut_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32438\,
            in1 => \N__36610\,
            in2 => \_gnd_net_\,
            in3 => \N__33258\,
            lcout => \Inst_core.n1705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i3_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001011010"
        )
    port map (
            in0 => \N__32396\,
            in1 => \N__32381\,
            in2 => \N__32360\,
            in3 => \N__33558\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37613\,
            ce => 'H',
            sr => \N__32255\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i9_4_lut_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32239\,
            in1 => \N__33010\,
            in2 => \N__32999\,
            in3 => \N__32977\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i15_4_lut_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32966\,
            in1 => \N__32798\,
            in2 => \N__32960\,
            in3 => \N__32864\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i11_4_lut_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32929\,
            in1 => \N__32908\,
            in2 => \N__32896\,
            in3 => \N__32875\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.i10_4_lut_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32854\,
            in1 => \N__32842\,
            in2 => \N__32830\,
            in3 => \N__32809\,
            lcout => \Inst_core.Inst_trigger.stages_1__Inst_stage.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__32792\,
            in1 => \N__32777\,
            in2 => \N__33302\,
            in3 => \N__32765\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0\,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7869\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__35099\,
            in1 => \N__33753\,
            in2 => \N__33338\,
            in3 => \N__32762\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7869\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7870\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__32759\,
            in1 => \N__32738\,
            in2 => \N__33780\,
            in3 => \N__32726\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7870\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7871\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i3_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__32723\,
            in1 => \N__33757\,
            in2 => \N__35123\,
            in3 => \N__32708\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7871\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7872\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__33224\,
            in1 => \N__33316\,
            in2 => \N__33781\,
            in3 => \N__33209\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7872\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7873\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__33206\,
            in1 => \N__33761\,
            in2 => \N__35143\,
            in3 => \N__33191\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7873\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7874\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__33188\,
            in1 => \N__33352\,
            in2 => \N__33782\,
            in3 => \N__33173\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7874\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7875\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__33170\,
            in1 => \N__33765\,
            in2 => \N__33152\,
            in3 => \N__33134\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7875\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7876\,
            clk => \N__37604\,
            ce => \N__33692\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i8_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__33131\,
            in1 => \N__33766\,
            in2 => \N__35171\,
            in3 => \N__33116\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7877\,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i9_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__33113\,
            in1 => \N__33098\,
            in2 => \N__33783\,
            in3 => \N__33086\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7877\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7878\,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i10_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__33083\,
            in1 => \N__33770\,
            in2 => \N__33065\,
            in3 => \N__33050\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7878\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7879\,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i11_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__33047\,
            in1 => \N__33029\,
            in2 => \N__33784\,
            in3 => \N__33017\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7879\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7880\,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i12_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__34283\,
            in1 => \N__33774\,
            in2 => \N__33863\,
            in3 => \N__33848\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7880\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7881\,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i13_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__33845\,
            in1 => \N__35156\,
            in2 => \N__33785\,
            in3 => \N__33824\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7881\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7882\,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i14_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__33821\,
            in1 => \N__33778\,
            in2 => \N__33803\,
            in3 => \N__33788\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7882\,
            carryout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n7883\,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i15_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__33779\,
            in1 => \N__33878\,
            in2 => \N__33710\,
            in3 => \N__33713\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37593\,
            ce => \N__33691\,
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011010100110"
        )
    port map (
            in0 => \N__33668\,
            in1 => \N__33647\,
            in2 => \N__33560\,
            in3 => \N__33467\,
            lcout => \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37579\,
            ce => 'H',
            sr => \N__33431\
        );

    \Inst_core.Inst_trigger.i3_4_lut_adj_78_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33419\,
            in1 => \N__33404\,
            in2 => \N__33392\,
            in3 => \N__33377\,
            lcout => \Inst_core.Inst_trigger.levelReg_1__N_590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i9_4_lut_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33353\,
            in1 => \N__33337\,
            in2 => \N__33320\,
            in3 => \N__33301\,
            lcout => OPEN,
            ltout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i15_4_lut_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33284\,
            in1 => \N__35105\,
            in2 => \N__33278\,
            in3 => \N__33275\,
            lcout => \Inst_core.n31_adj_1132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.i10_4_lut_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35167\,
            in1 => \N__35155\,
            in2 => \N__35144\,
            in3 => \N__35122\,
            lcout => \Inst_core.Inst_trigger.stages_0__Inst_stage.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i2_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34261\,
            in1 => \_gnd_net_\,
            in2 => \N__34124\,
            in3 => \N__35095\,
            lcout => \configRegister_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i17_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36160\,
            in1 => \N__34115\,
            in2 => \_gnd_net_\,
            in3 => \N__35083\,
            lcout => \configRegister_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_eia232.Inst_receiver.dataBuf_i12_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__34568\,
            in1 => \N__34964\,
            in2 => \N__34850\,
            in3 => \N__35312\,
            lcout => cmd_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i6_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34520\,
            in1 => \N__34432\,
            in2 => \_gnd_net_\,
            in3 => \N__34294\,
            lcout => \valueRegister_6_adj_1290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i13_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34113\,
            in1 => \N__35311\,
            in2 => \_gnd_net_\,
            in3 => \N__34279\,
            lcout => \configRegister_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i1_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35505\,
            in1 => \N__34260\,
            in2 => \_gnd_net_\,
            in3 => \N__34138\,
            lcout => bwd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i16_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34114\,
            in1 => \N__33940\,
            in2 => \_gnd_net_\,
            in3 => \N__33874\,
            lcout => \configRegister_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i17_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36161\,
            in1 => \N__35849\,
            in2 => \_gnd_net_\,
            in3 => \N__36118\,
            lcout => \configRegister_16_adj_1344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i0_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36091\,
            in1 => \N__35995\,
            in2 => \_gnd_net_\,
            in3 => \N__36010\,
            lcout => \valueRegister_0_adj_1376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35442\,
            in1 => \N__35996\,
            in2 => \_gnd_net_\,
            in3 => \N__35872\,
            lcout => bwd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i24_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35539\,
            in1 => \N__35848\,
            in2 => \_gnd_net_\,
            in3 => \N__35681\,
            lcout => \configRegister_26_adj_1337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.bwd_i0_i12_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35443\,
            in1 => \N__35309\,
            in2 => \_gnd_net_\,
            in3 => \N__35233\,
            lcout => bwd_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.state_FSM_i2_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__36450\,
            in1 => \N__36705\,
            in2 => \N__36716\,
            in3 => \N__36689\,
            lcout => send,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37603\,
            ce => 'H',
            sr => \N__36875\
        );

    \Inst_core.Inst_controller.state_FSM_i1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__36688\,
            in1 => \N__35197\,
            in2 => \N__36707\,
            in3 => \N__35219\,
            lcout => \Inst_core.Inst_controller.n320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37603\,
            ce => 'H',
            sr => \N__36875\
        );

    \Inst_core.Inst_controller.state_FSM_i0_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__36321\,
            in1 => \N__35215\,
            in2 => \N__35198\,
            in3 => \N__35185\,
            lcout => \Inst_core.Inst_controller.n321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37603\,
            ce => 'H',
            sr => \N__36875\
        );

    \Inst_core.Inst_controller.state_FSM_i3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110010100000"
        )
    port map (
            in0 => \N__35186\,
            in1 => \N__36731\,
            in2 => \N__36339\,
            in3 => \N__36451\,
            lcout => \Inst_core.n318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37603\,
            ce => 'H',
            sr => \N__36875\
        );

    \Inst_core.Inst_controller.i1605_3_lut_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__36452\,
            in1 => \N__36325\,
            in2 => \_gnd_net_\,
            in3 => \N__36706\,
            lcout => debugleds_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i5479_2_lut_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36730\,
            in2 => \_gnd_net_\,
            in3 => \N__36320\,
            lcout => \Inst_core.Inst_controller.nstate_1_N_825_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i1608_2_lut_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36701\,
            in2 => \_gnd_net_\,
            in3 => \N__36687\,
            lcout => \Inst_core.Inst_controller.n2717\,
            ltout => \Inst_core.Inst_controller.n2717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.i5504_3_lut_4_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__36557\,
            in1 => \N__36449\,
            in2 => \N__36428\,
            in3 => \N__36319\,
            lcout => \Inst_core.Inst_controller.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Inst_core.Inst_controller.counter__i0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36275\,
            in2 => \_gnd_net_\,
            in3 => \N__36260\,
            lcout => \Inst_core.Inst_controller.counter_0\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \Inst_core.Inst_controller.n7845\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36257\,
            in2 => \_gnd_net_\,
            in3 => \N__36239\,
            lcout => \Inst_core.Inst_controller.counter_1\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7845\,
            carryout => \Inst_core.Inst_controller.n7846\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36236\,
            in2 => \_gnd_net_\,
            in3 => \N__36218\,
            lcout => \Inst_core.Inst_controller.counter_2\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7846\,
            carryout => \Inst_core.Inst_controller.n7847\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36204\,
            in2 => \_gnd_net_\,
            in3 => \N__36188\,
            lcout => \Inst_core.Inst_controller.counter_3\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7847\,
            carryout => \Inst_core.Inst_controller.n7848\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i4_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37100\,
            in2 => \_gnd_net_\,
            in3 => \N__37082\,
            lcout => \Inst_core.Inst_controller.counter_4\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7848\,
            carryout => \Inst_core.Inst_controller.n7849\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i5_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37071\,
            in2 => \_gnd_net_\,
            in3 => \N__37055\,
            lcout => \Inst_core.Inst_controller.counter_5\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7849\,
            carryout => \Inst_core.Inst_controller.n7850\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i6_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37044\,
            in2 => \_gnd_net_\,
            in3 => \N__37028\,
            lcout => \Inst_core.Inst_controller.counter_6\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7850\,
            carryout => \Inst_core.Inst_controller.n7851\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i7_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37014\,
            in2 => \_gnd_net_\,
            in3 => \N__36992\,
            lcout => \Inst_core.Inst_controller.counter_7\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7851\,
            carryout => \Inst_core.Inst_controller.n7852\,
            clk => \N__37612\,
            ce => \N__37157\,
            sr => \N__37116\
        );

    \Inst_core.Inst_controller.counter__i8_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36978\,
            in2 => \_gnd_net_\,
            in3 => \N__36956\,
            lcout => \Inst_core.Inst_controller.counter_8\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \Inst_core.Inst_controller.n7853\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i9_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36946\,
            in2 => \_gnd_net_\,
            in3 => \N__36932\,
            lcout => \Inst_core.Inst_controller.counter_9\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7853\,
            carryout => \Inst_core.Inst_controller.n7854\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i10_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36921\,
            in2 => \_gnd_net_\,
            in3 => \N__36905\,
            lcout => \Inst_core.Inst_controller.counter_10\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7854\,
            carryout => \Inst_core.Inst_controller.n7855\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i11_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36894\,
            in2 => \_gnd_net_\,
            in3 => \N__36878\,
            lcout => \Inst_core.Inst_controller.counter_11\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7855\,
            carryout => \Inst_core.Inst_controller.n7856\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i12_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37789\,
            in2 => \_gnd_net_\,
            in3 => \N__37775\,
            lcout => \Inst_core.Inst_controller.counter_12\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7856\,
            carryout => \Inst_core.Inst_controller.n7857\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i13_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37765\,
            in2 => \_gnd_net_\,
            in3 => \N__37751\,
            lcout => \Inst_core.Inst_controller.counter_13\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7857\,
            carryout => \Inst_core.Inst_controller.n7858\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i14_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37741\,
            in2 => \_gnd_net_\,
            in3 => \N__37727\,
            lcout => \Inst_core.Inst_controller.counter_14\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7858\,
            carryout => \Inst_core.Inst_controller.n7859\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i15_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37719\,
            in2 => \_gnd_net_\,
            in3 => \N__37700\,
            lcout => \Inst_core.Inst_controller.counter_15\,
            ltout => OPEN,
            carryin => \Inst_core.Inst_controller.n7859\,
            carryout => \Inst_core.Inst_controller.n7860\,
            clk => \N__37619\,
            ce => \N__37156\,
            sr => \N__37117\
        );

    \Inst_core.Inst_controller.counter__i16_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37686\,
            in2 => \_gnd_net_\,
            in3 => \N__37670\,
            lcout => \Inst_core.Inst_controller.counter_16\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \Inst_core.Inst_controller.n7861\,
            clk => \N__37625\,
            ce => \N__37152\,
            sr => \N__37124\
        );

    \Inst_core.Inst_controller.counter__i17_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37656\,
            in2 => \_gnd_net_\,
            in3 => \N__37667\,
            lcout => \Inst_core.Inst_controller.counter_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37625\,
            ce => \N__37152\,
            sr => \N__37124\
        );
end \INTERFACE\;
