// ******************************************************************************

// iCEcube Netlister

// Version:            2016.02.27810

// Build Date:         Jan 29 2016 01:59:28

// File Generated:     Aug 24 2016 00:01:55

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "la" view "INTERFACE"

module la (
    debugleds,
    testcnt,
    \input ,
    xtalClock,
    tx,
    rx,
    ready50,
    exClock);

    output [1:0] debugleds;
    output [7:0] testcnt;
    input [7:0] input;
    input xtalClock;
    output tx;
    input rx;
    output ready50;
    input exClock;

    wire N__38006;
    wire N__38005;
    wire N__38004;
    wire N__37995;
    wire N__37994;
    wire N__37993;
    wire N__37986;
    wire N__37985;
    wire N__37984;
    wire N__37977;
    wire N__37976;
    wire N__37975;
    wire N__37968;
    wire N__37967;
    wire N__37966;
    wire N__37959;
    wire N__37958;
    wire N__37957;
    wire N__37950;
    wire N__37949;
    wire N__37948;
    wire N__37941;
    wire N__37940;
    wire N__37939;
    wire N__37932;
    wire N__37931;
    wire N__37930;
    wire N__37923;
    wire N__37922;
    wire N__37921;
    wire N__37914;
    wire N__37913;
    wire N__37912;
    wire N__37905;
    wire N__37904;
    wire N__37903;
    wire N__37896;
    wire N__37895;
    wire N__37894;
    wire N__37887;
    wire N__37886;
    wire N__37885;
    wire N__37878;
    wire N__37877;
    wire N__37876;
    wire N__37869;
    wire N__37868;
    wire N__37867;
    wire N__37860;
    wire N__37859;
    wire N__37858;
    wire N__37851;
    wire N__37850;
    wire N__37849;
    wire N__37842;
    wire N__37841;
    wire N__37840;
    wire N__37833;
    wire N__37832;
    wire N__37831;
    wire N__37824;
    wire N__37823;
    wire N__37822;
    wire N__37815;
    wire N__37814;
    wire N__37813;
    wire N__37796;
    wire N__37795;
    wire N__37790;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37775;
    wire N__37772;
    wire N__37771;
    wire N__37766;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37751;
    wire N__37748;
    wire N__37747;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37727;
    wire N__37724;
    wire N__37723;
    wire N__37720;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37705;
    wire N__37700;
    wire N__37697;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37686;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37636;
    wire N__37633;
    wire N__37628;
    wire N__37627;
    wire N__37626;
    wire N__37625;
    wire N__37624;
    wire N__37623;
    wire N__37622;
    wire N__37621;
    wire N__37620;
    wire N__37619;
    wire N__37618;
    wire N__37617;
    wire N__37616;
    wire N__37615;
    wire N__37614;
    wire N__37613;
    wire N__37612;
    wire N__37611;
    wire N__37610;
    wire N__37609;
    wire N__37608;
    wire N__37607;
    wire N__37606;
    wire N__37605;
    wire N__37604;
    wire N__37603;
    wire N__37602;
    wire N__37601;
    wire N__37600;
    wire N__37599;
    wire N__37598;
    wire N__37597;
    wire N__37596;
    wire N__37595;
    wire N__37594;
    wire N__37593;
    wire N__37592;
    wire N__37591;
    wire N__37590;
    wire N__37589;
    wire N__37588;
    wire N__37587;
    wire N__37586;
    wire N__37585;
    wire N__37584;
    wire N__37583;
    wire N__37582;
    wire N__37581;
    wire N__37580;
    wire N__37579;
    wire N__37578;
    wire N__37577;
    wire N__37576;
    wire N__37575;
    wire N__37574;
    wire N__37573;
    wire N__37572;
    wire N__37571;
    wire N__37570;
    wire N__37569;
    wire N__37568;
    wire N__37567;
    wire N__37566;
    wire N__37565;
    wire N__37564;
    wire N__37563;
    wire N__37562;
    wire N__37561;
    wire N__37560;
    wire N__37559;
    wire N__37558;
    wire N__37557;
    wire N__37556;
    wire N__37555;
    wire N__37554;
    wire N__37553;
    wire N__37552;
    wire N__37551;
    wire N__37550;
    wire N__37549;
    wire N__37548;
    wire N__37547;
    wire N__37546;
    wire N__37545;
    wire N__37544;
    wire N__37543;
    wire N__37542;
    wire N__37541;
    wire N__37540;
    wire N__37539;
    wire N__37538;
    wire N__37537;
    wire N__37536;
    wire N__37535;
    wire N__37534;
    wire N__37533;
    wire N__37532;
    wire N__37531;
    wire N__37530;
    wire N__37529;
    wire N__37528;
    wire N__37527;
    wire N__37526;
    wire N__37525;
    wire N__37524;
    wire N__37523;
    wire N__37522;
    wire N__37521;
    wire N__37520;
    wire N__37519;
    wire N__37518;
    wire N__37517;
    wire N__37516;
    wire N__37515;
    wire N__37514;
    wire N__37513;
    wire N__37512;
    wire N__37511;
    wire N__37510;
    wire N__37509;
    wire N__37508;
    wire N__37507;
    wire N__37506;
    wire N__37505;
    wire N__37504;
    wire N__37503;
    wire N__37502;
    wire N__37501;
    wire N__37500;
    wire N__37499;
    wire N__37498;
    wire N__37497;
    wire N__37496;
    wire N__37495;
    wire N__37494;
    wire N__37493;
    wire N__37492;
    wire N__37491;
    wire N__37490;
    wire N__37489;
    wire N__37488;
    wire N__37487;
    wire N__37486;
    wire N__37485;
    wire N__37484;
    wire N__37483;
    wire N__37482;
    wire N__37481;
    wire N__37480;
    wire N__37479;
    wire N__37478;
    wire N__37477;
    wire N__37476;
    wire N__37475;
    wire N__37474;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37156;
    wire N__37153;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37135;
    wire N__37132;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37117;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37100;
    wire N__37099;
    wire N__37098;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37082;
    wire N__37079;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37071;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37055;
    wire N__37052;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37044;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37028;
    wire N__37025;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36992;
    wire N__36989;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36956;
    wire N__36953;
    wire N__36952;
    wire N__36947;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36932;
    wire N__36929;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36921;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36905;
    wire N__36902;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36894;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36878;
    wire N__36875;
    wire N__36874;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36864;
    wire N__36861;
    wire N__36860;
    wire N__36859;
    wire N__36858;
    wire N__36855;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36823;
    wire N__36818;
    wire N__36813;
    wire N__36812;
    wire N__36809;
    wire N__36808;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36746;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36730;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36706;
    wire N__36705;
    wire N__36702;
    wire N__36701;
    wire N__36692;
    wire N__36689;
    wire N__36688;
    wire N__36687;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36664;
    wire N__36663;
    wire N__36662;
    wire N__36659;
    wire N__36658;
    wire N__36657;
    wire N__36656;
    wire N__36651;
    wire N__36648;
    wire N__36647;
    wire N__36646;
    wire N__36645;
    wire N__36644;
    wire N__36643;
    wire N__36640;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36634;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36626;
    wire N__36625;
    wire N__36622;
    wire N__36613;
    wire N__36612;
    wire N__36611;
    wire N__36610;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36598;
    wire N__36589;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36566;
    wire N__36565;
    wire N__36564;
    wire N__36563;
    wire N__36562;
    wire N__36561;
    wire N__36558;
    wire N__36557;
    wire N__36554;
    wire N__36553;
    wire N__36548;
    wire N__36543;
    wire N__36534;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36512;
    wire N__36509;
    wire N__36508;
    wire N__36503;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36479;
    wire N__36474;
    wire N__36469;
    wire N__36462;
    wire N__36459;
    wire N__36452;
    wire N__36451;
    wire N__36450;
    wire N__36449;
    wire N__36448;
    wire N__36447;
    wire N__36438;
    wire N__36433;
    wire N__36428;
    wire N__36425;
    wire N__36424;
    wire N__36423;
    wire N__36422;
    wire N__36415;
    wire N__36414;
    wire N__36413;
    wire N__36412;
    wire N__36411;
    wire N__36410;
    wire N__36409;
    wire N__36408;
    wire N__36407;
    wire N__36406;
    wire N__36403;
    wire N__36402;
    wire N__36401;
    wire N__36400;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36375;
    wire N__36370;
    wire N__36363;
    wire N__36358;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36339;
    wire N__36334;
    wire N__36331;
    wire N__36326;
    wire N__36325;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36318;
    wire N__36317;
    wire N__36310;
    wire N__36305;
    wire N__36298;
    wire N__36293;
    wire N__36290;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36274;
    wire N__36273;
    wire N__36270;
    wire N__36265;
    wire N__36260;
    wire N__36257;
    wire N__36256;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36204;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36188;
    wire N__36185;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36177;
    wire N__36176;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36162;
    wire N__36161;
    wire N__36160;
    wire N__36155;
    wire N__36152;
    wire N__36147;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36104;
    wire N__36103;
    wire N__36100;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36092;
    wire N__36091;
    wire N__36090;
    wire N__36089;
    wire N__36088;
    wire N__36085;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36057;
    wire N__36052;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__35999;
    wire N__35998;
    wire N__35997;
    wire N__35996;
    wire N__35995;
    wire N__35990;
    wire N__35989;
    wire N__35988;
    wire N__35985;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35958;
    wire N__35957;
    wire N__35956;
    wire N__35955;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35929;
    wire N__35928;
    wire N__35927;
    wire N__35926;
    wire N__35925;
    wire N__35922;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35904;
    wire N__35901;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35873;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35858;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35854;
    wire N__35853;
    wire N__35852;
    wire N__35851;
    wire N__35850;
    wire N__35849;
    wire N__35848;
    wire N__35845;
    wire N__35836;
    wire N__35835;
    wire N__35834;
    wire N__35833;
    wire N__35832;
    wire N__35831;
    wire N__35826;
    wire N__35821;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35813;
    wire N__35808;
    wire N__35803;
    wire N__35802;
    wire N__35801;
    wire N__35800;
    wire N__35799;
    wire N__35796;
    wire N__35795;
    wire N__35794;
    wire N__35791;
    wire N__35790;
    wire N__35787;
    wire N__35782;
    wire N__35779;
    wire N__35774;
    wire N__35771;
    wire N__35766;
    wire N__35763;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35733;
    wire N__35730;
    wire N__35725;
    wire N__35720;
    wire N__35715;
    wire N__35708;
    wire N__35701;
    wire N__35698;
    wire N__35691;
    wire N__35688;
    wire N__35681;
    wire N__35680;
    wire N__35677;
    wire N__35676;
    wire N__35673;
    wire N__35672;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35651;
    wire N__35644;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35612;
    wire N__35611;
    wire N__35610;
    wire N__35607;
    wire N__35606;
    wire N__35605;
    wire N__35602;
    wire N__35601;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35578;
    wire N__35575;
    wire N__35570;
    wire N__35567;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35548;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35536;
    wire N__35529;
    wire N__35526;
    wire N__35519;
    wire N__35518;
    wire N__35517;
    wire N__35516;
    wire N__35515;
    wire N__35514;
    wire N__35513;
    wire N__35512;
    wire N__35511;
    wire N__35510;
    wire N__35509;
    wire N__35508;
    wire N__35507;
    wire N__35506;
    wire N__35505;
    wire N__35500;
    wire N__35497;
    wire N__35492;
    wire N__35479;
    wire N__35478;
    wire N__35477;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35466;
    wire N__35465;
    wire N__35462;
    wire N__35453;
    wire N__35448;
    wire N__35445;
    wire N__35444;
    wire N__35443;
    wire N__35442;
    wire N__35441;
    wire N__35434;
    wire N__35433;
    wire N__35432;
    wire N__35427;
    wire N__35422;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35383;
    wire N__35378;
    wire N__35375;
    wire N__35366;
    wire N__35365;
    wire N__35364;
    wire N__35357;
    wire N__35354;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35307;
    wire N__35302;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35290;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35254;
    wire N__35251;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35219;
    wire N__35216;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35197;
    wire N__35194;
    wire N__35189;
    wire N__35186;
    wire N__35185;
    wire N__35184;
    wire N__35179;
    wire N__35176;
    wire N__35171;
    wire N__35168;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35156;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35144;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35123;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35096;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35084;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35069;
    wire N__35068;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35060;
    wire N__35059;
    wire N__35058;
    wire N__35057;
    wire N__35056;
    wire N__35055;
    wire N__35054;
    wire N__35053;
    wire N__35052;
    wire N__35051;
    wire N__35050;
    wire N__35049;
    wire N__35048;
    wire N__35047;
    wire N__35046;
    wire N__35045;
    wire N__35042;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35026;
    wire N__35023;
    wire N__35018;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35006;
    wire N__34997;
    wire N__34996;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34966;
    wire N__34965;
    wire N__34964;
    wire N__34963;
    wire N__34962;
    wire N__34961;
    wire N__34960;
    wire N__34959;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34936;
    wire N__34935;
    wire N__34934;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34911;
    wire N__34906;
    wire N__34901;
    wire N__34898;
    wire N__34891;
    wire N__34886;
    wire N__34881;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34857;
    wire N__34850;
    wire N__34847;
    wire N__34846;
    wire N__34845;
    wire N__34844;
    wire N__34843;
    wire N__34842;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34836;
    wire N__34827;
    wire N__34826;
    wire N__34825;
    wire N__34822;
    wire N__34821;
    wire N__34820;
    wire N__34819;
    wire N__34818;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34810;
    wire N__34809;
    wire N__34806;
    wire N__34805;
    wire N__34804;
    wire N__34803;
    wire N__34802;
    wire N__34801;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34778;
    wire N__34777;
    wire N__34776;
    wire N__34775;
    wire N__34774;
    wire N__34773;
    wire N__34768;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34747;
    wire N__34744;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34725;
    wire N__34722;
    wire N__34717;
    wire N__34712;
    wire N__34707;
    wire N__34706;
    wire N__34703;
    wire N__34702;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34687;
    wire N__34680;
    wire N__34675;
    wire N__34672;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34642;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34622;
    wire N__34615;
    wire N__34612;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34592;
    wire N__34591;
    wire N__34588;
    wire N__34583;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34524;
    wire N__34523;
    wire N__34522;
    wire N__34521;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34451;
    wire N__34448;
    wire N__34443;
    wire N__34440;
    wire N__34433;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34422;
    wire N__34421;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34410;
    wire N__34409;
    wire N__34408;
    wire N__34405;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34376;
    wire N__34373;
    wire N__34368;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34356;
    wire N__34353;
    wire N__34348;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34327;
    wire N__34324;
    wire N__34317;
    wire N__34308;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34283;
    wire N__34280;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34268;
    wire N__34267;
    wire N__34266;
    wire N__34263;
    wire N__34262;
    wire N__34261;
    wire N__34260;
    wire N__34259;
    wire N__34258;
    wire N__34257;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34241;
    wire N__34238;
    wire N__34237;
    wire N__34232;
    wire N__34231;
    wire N__34228;
    wire N__34227;
    wire N__34226;
    wire N__34223;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34206;
    wire N__34205;
    wire N__34202;
    wire N__34197;
    wire N__34196;
    wire N__34191;
    wire N__34188;
    wire N__34183;
    wire N__34180;
    wire N__34179;
    wire N__34176;
    wire N__34171;
    wire N__34168;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34142;
    wire N__34139;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34124;
    wire N__34123;
    wire N__34122;
    wire N__34121;
    wire N__34120;
    wire N__34119;
    wire N__34116;
    wire N__34115;
    wire N__34114;
    wire N__34113;
    wire N__34108;
    wire N__34107;
    wire N__34106;
    wire N__34105;
    wire N__34104;
    wire N__34103;
    wire N__34102;
    wire N__34101;
    wire N__34100;
    wire N__34099;
    wire N__34098;
    wire N__34097;
    wire N__34096;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34085;
    wire N__34084;
    wire N__34075;
    wire N__34072;
    wire N__34067;
    wire N__34064;
    wire N__34057;
    wire N__34050;
    wire N__34047;
    wire N__34046;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34015;
    wire N__34012;
    wire N__34007;
    wire N__34002;
    wire N__33999;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33961;
    wire N__33956;
    wire N__33951;
    wire N__33948;
    wire N__33941;
    wire N__33940;
    wire N__33937;
    wire N__33936;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33928;
    wire N__33923;
    wire N__33918;
    wire N__33915;
    wire N__33914;
    wire N__33913;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33898;
    wire N__33893;
    wire N__33888;
    wire N__33885;
    wire N__33878;
    wire N__33875;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33863;
    wire N__33860;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33803;
    wire N__33800;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33788;
    wire N__33785;
    wire N__33784;
    wire N__33783;
    wire N__33782;
    wire N__33781;
    wire N__33780;
    wire N__33779;
    wire N__33778;
    wire N__33775;
    wire N__33774;
    wire N__33771;
    wire N__33770;
    wire N__33767;
    wire N__33766;
    wire N__33765;
    wire N__33762;
    wire N__33761;
    wire N__33758;
    wire N__33757;
    wire N__33754;
    wire N__33753;
    wire N__33736;
    wire N__33721;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33692;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33668;
    wire N__33665;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33653;
    wire N__33652;
    wire N__33651;
    wire N__33648;
    wire N__33647;
    wire N__33646;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33638;
    wire N__33635;
    wire N__33634;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33585;
    wire N__33582;
    wire N__33577;
    wire N__33574;
    wire N__33569;
    wire N__33560;
    wire N__33559;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33553;
    wire N__33552;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33481;
    wire N__33478;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33453;
    wire N__33448;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33364;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33338;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33320;
    wire N__33317;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33302;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33266;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33258;
    wire N__33253;
    wire N__33250;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33224;
    wire N__33221;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33152;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33134;
    wire N__33131;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33098;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33065;
    wire N__33062;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33041;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33029;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__32999;
    wire N__32996;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32981;
    wire N__32978;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32950;
    wire N__32949;
    wire N__32948;
    wire N__32947;
    wire N__32944;
    wire N__32935;
    wire N__32930;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32912;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32897;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32887;
    wire N__32884;
    wire N__32879;
    wire N__32876;
    wire N__32875;
    wire N__32872;
    wire N__32869;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32854;
    wire N__32851;
    wire N__32848;
    wire N__32843;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32813;
    wire N__32810;
    wire N__32809;
    wire N__32806;
    wire N__32803;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32738;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32719;
    wire N__32716;
    wire N__32713;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32662;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32621;
    wire N__32620;
    wire N__32613;
    wire N__32610;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32542;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32524;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32489;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32477;
    wire N__32474;
    wire N__32473;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32450;
    wire N__32449;
    wire N__32444;
    wire N__32441;
    wire N__32440;
    wire N__32439;
    wire N__32438;
    wire N__32435;
    wire N__32434;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32416;
    wire N__32413;
    wire N__32408;
    wire N__32405;
    wire N__32396;
    wire N__32393;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32374;
    wire N__32373;
    wire N__32370;
    wire N__32365;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32353;
    wire N__32352;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32344;
    wire N__32343;
    wire N__32340;
    wire N__32339;
    wire N__32338;
    wire N__32337;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32313;
    wire N__32310;
    wire N__32305;
    wire N__32300;
    wire N__32297;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32275;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32213;
    wire N__32210;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32198;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32190;
    wire N__32187;
    wire N__32182;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32101;
    wire N__32098;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32081;
    wire N__32080;
    wire N__32077;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32060;
    wire N__32057;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32032;
    wire N__32027;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31963;
    wire N__31962;
    wire N__31961;
    wire N__31960;
    wire N__31957;
    wire N__31956;
    wire N__31955;
    wire N__31954;
    wire N__31953;
    wire N__31950;
    wire N__31949;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31904;
    wire N__31897;
    wire N__31896;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31884;
    wire N__31881;
    wire N__31876;
    wire N__31873;
    wire N__31862;
    wire N__31861;
    wire N__31858;
    wire N__31857;
    wire N__31854;
    wire N__31849;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31805;
    wire N__31804;
    wire N__31801;
    wire N__31800;
    wire N__31797;
    wire N__31796;
    wire N__31795;
    wire N__31794;
    wire N__31791;
    wire N__31790;
    wire N__31789;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31729;
    wire N__31726;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31701;
    wire N__31698;
    wire N__31693;
    wire N__31688;
    wire N__31687;
    wire N__31684;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31663;
    wire N__31660;
    wire N__31655;
    wire N__31654;
    wire N__31651;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31618;
    wire N__31617;
    wire N__31614;
    wire N__31609;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31553;
    wire N__31550;
    wire N__31549;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31529;
    wire N__31528;
    wire N__31525;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31510;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31483;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31436;
    wire N__31435;
    wire N__31432;
    wire N__31429;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31406;
    wire N__31403;
    wire N__31402;
    wire N__31399;
    wire N__31398;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31387;
    wire N__31384;
    wire N__31383;
    wire N__31380;
    wire N__31375;
    wire N__31374;
    wire N__31371;
    wire N__31370;
    wire N__31369;
    wire N__31368;
    wire N__31365;
    wire N__31364;
    wire N__31361;
    wire N__31356;
    wire N__31353;
    wire N__31352;
    wire N__31351;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31332;
    wire N__31325;
    wire N__31324;
    wire N__31323;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31311;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31275;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31251;
    wire N__31248;
    wire N__31243;
    wire N__31232;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31202;
    wire N__31199;
    wire N__31198;
    wire N__31197;
    wire N__31196;
    wire N__31193;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31185;
    wire N__31182;
    wire N__31177;
    wire N__31172;
    wire N__31169;
    wire N__31168;
    wire N__31167;
    wire N__31166;
    wire N__31165;
    wire N__31164;
    wire N__31163;
    wire N__31158;
    wire N__31153;
    wire N__31146;
    wire N__31141;
    wire N__31140;
    wire N__31139;
    wire N__31138;
    wire N__31137;
    wire N__31136;
    wire N__31133;
    wire N__31124;
    wire N__31115;
    wire N__31114;
    wire N__31113;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31107;
    wire N__31106;
    wire N__31105;
    wire N__31104;
    wire N__31103;
    wire N__31102;
    wire N__31099;
    wire N__31094;
    wire N__31093;
    wire N__31092;
    wire N__31091;
    wire N__31090;
    wire N__31089;
    wire N__31082;
    wire N__31077;
    wire N__31072;
    wire N__31067;
    wire N__31062;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31043;
    wire N__31040;
    wire N__31035;
    wire N__31032;
    wire N__31031;
    wire N__31028;
    wire N__31023;
    wire N__31016;
    wire N__31013;
    wire N__31008;
    wire N__31005;
    wire N__30998;
    wire N__30993;
    wire N__30992;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30940;
    wire N__30937;
    wire N__30936;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30928;
    wire N__30925;
    wire N__30924;
    wire N__30923;
    wire N__30922;
    wire N__30921;
    wire N__30918;
    wire N__30913;
    wire N__30910;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30875;
    wire N__30872;
    wire N__30867;
    wire N__30864;
    wire N__30859;
    wire N__30854;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30827;
    wire N__30824;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30816;
    wire N__30813;
    wire N__30808;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30749;
    wire N__30746;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30731;
    wire N__30728;
    wire N__30727;
    wire N__30722;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30707;
    wire N__30704;
    wire N__30703;
    wire N__30700;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30670;
    wire N__30667;
    wire N__30666;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30637;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30622;
    wire N__30617;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30595;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30583;
    wire N__30580;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30557;
    wire N__30556;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30541;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30523;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30508;
    wire N__30503;
    wire N__30502;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30487;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30467;
    wire N__30466;
    wire N__30463;
    wire N__30462;
    wire N__30461;
    wire N__30458;
    wire N__30457;
    wire N__30456;
    wire N__30453;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30409;
    wire N__30406;
    wire N__30405;
    wire N__30402;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30373;
    wire N__30366;
    wire N__30359;
    wire N__30358;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30347;
    wire N__30346;
    wire N__30345;
    wire N__30344;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30297;
    wire N__30296;
    wire N__30293;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30268;
    wire N__30263;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30191;
    wire N__30188;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30115;
    wire N__30114;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30100;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30069;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30035;
    wire N__30034;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30012;
    wire N__30009;
    wire N__30002;
    wire N__30001;
    wire N__29998;
    wire N__29993;
    wire N__29990;
    wire N__29989;
    wire N__29988;
    wire N__29985;
    wire N__29980;
    wire N__29975;
    wire N__29972;
    wire N__29971;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29936;
    wire N__29933;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29918;
    wire N__29915;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29813;
    wire N__29810;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29802;
    wire N__29799;
    wire N__29794;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29765;
    wire N__29764;
    wire N__29759;
    wire N__29758;
    wire N__29757;
    wire N__29756;
    wire N__29753;
    wire N__29752;
    wire N__29751;
    wire N__29746;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29725;
    wire N__29714;
    wire N__29713;
    wire N__29712;
    wire N__29711;
    wire N__29708;
    wire N__29707;
    wire N__29706;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29680;
    wire N__29679;
    wire N__29678;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29672;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29626;
    wire N__29625;
    wire N__29624;
    wire N__29623;
    wire N__29616;
    wire N__29611;
    wire N__29606;
    wire N__29603;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29584;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29555;
    wire N__29554;
    wire N__29549;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29541;
    wire N__29540;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29528;
    wire N__29527;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29502;
    wire N__29495;
    wire N__29494;
    wire N__29491;
    wire N__29490;
    wire N__29489;
    wire N__29484;
    wire N__29483;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29475;
    wire N__29472;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29457;
    wire N__29452;
    wire N__29449;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29414;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29399;
    wire N__29396;
    wire N__29395;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29384;
    wire N__29383;
    wire N__29382;
    wire N__29379;
    wire N__29374;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29356;
    wire N__29355;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29333;
    wire N__29332;
    wire N__29331;
    wire N__29330;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29324;
    wire N__29321;
    wire N__29320;
    wire N__29319;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29311;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29300;
    wire N__29299;
    wire N__29296;
    wire N__29295;
    wire N__29294;
    wire N__29293;
    wire N__29292;
    wire N__29291;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29279;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29267;
    wire N__29262;
    wire N__29259;
    wire N__29254;
    wire N__29253;
    wire N__29252;
    wire N__29251;
    wire N__29250;
    wire N__29243;
    wire N__29240;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29224;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29206;
    wire N__29197;
    wire N__29194;
    wire N__29187;
    wire N__29184;
    wire N__29179;
    wire N__29176;
    wire N__29171;
    wire N__29164;
    wire N__29159;
    wire N__29152;
    wire N__29147;
    wire N__29144;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29132;
    wire N__29131;
    wire N__29130;
    wire N__29129;
    wire N__29128;
    wire N__29127;
    wire N__29124;
    wire N__29123;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29115;
    wire N__29114;
    wire N__29111;
    wire N__29110;
    wire N__29109;
    wire N__29108;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29097;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29064;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29044;
    wire N__29041;
    wire N__29036;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29007;
    wire N__29000;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28964;
    wire N__28963;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28955;
    wire N__28954;
    wire N__28951;
    wire N__28946;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28928;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28913;
    wire N__28912;
    wire N__28911;
    wire N__28910;
    wire N__28909;
    wire N__28904;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28885;
    wire N__28880;
    wire N__28879;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28793;
    wire N__28790;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28772;
    wire N__28769;
    wire N__28768;
    wire N__28767;
    wire N__28766;
    wire N__28763;
    wire N__28762;
    wire N__28761;
    wire N__28758;
    wire N__28757;
    wire N__28754;
    wire N__28753;
    wire N__28750;
    wire N__28749;
    wire N__28746;
    wire N__28745;
    wire N__28744;
    wire N__28743;
    wire N__28726;
    wire N__28723;
    wire N__28722;
    wire N__28719;
    wire N__28718;
    wire N__28715;
    wire N__28714;
    wire N__28711;
    wire N__28710;
    wire N__28705;
    wire N__28690;
    wire N__28687;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28661;
    wire N__28658;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28646;
    wire N__28643;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28635;
    wire N__28632;
    wire N__28627;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28553;
    wire N__28550;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28406;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28394;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28340;
    wire N__28339;
    wire N__28338;
    wire N__28337;
    wire N__28334;
    wire N__28327;
    wire N__28326;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28310;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28259;
    wire N__28256;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28192;
    wire N__28191;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28179;
    wire N__28178;
    wire N__28177;
    wire N__28176;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28136;
    wire N__28133;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28121;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28113;
    wire N__28110;
    wire N__28105;
    wire N__28102;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28087;
    wire N__28086;
    wire N__28085;
    wire N__28082;
    wire N__28081;
    wire N__28078;
    wire N__28077;
    wire N__28076;
    wire N__28073;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28029;
    wire N__28028;
    wire N__28027;
    wire N__28024;
    wire N__28019;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27880;
    wire N__27877;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27850;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27827;
    wire N__27824;
    wire N__27823;
    wire N__27822;
    wire N__27819;
    wire N__27814;
    wire N__27809;
    wire N__27806;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27756;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27724;
    wire N__27723;
    wire N__27720;
    wire N__27715;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27700;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27680;
    wire N__27677;
    wire N__27676;
    wire N__27675;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27649;
    wire N__27648;
    wire N__27645;
    wire N__27640;
    wire N__27635;
    wire N__27632;
    wire N__27631;
    wire N__27630;
    wire N__27627;
    wire N__27622;
    wire N__27617;
    wire N__27614;
    wire N__27613;
    wire N__27612;
    wire N__27609;
    wire N__27604;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27592;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27553;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27526;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27502;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27479;
    wire N__27476;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27437;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27361;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27340;
    wire N__27337;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27316;
    wire N__27315;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27299;
    wire N__27296;
    wire N__27295;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27280;
    wire N__27275;
    wire N__27274;
    wire N__27271;
    wire N__27266;
    wire N__27263;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27248;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27208;
    wire N__27207;
    wire N__27206;
    wire N__27205;
    wire N__27202;
    wire N__27201;
    wire N__27200;
    wire N__27199;
    wire N__27198;
    wire N__27197;
    wire N__27194;
    wire N__27193;
    wire N__27192;
    wire N__27191;
    wire N__27188;
    wire N__27183;
    wire N__27180;
    wire N__27175;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27143;
    wire N__27142;
    wire N__27141;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27129;
    wire N__27124;
    wire N__27121;
    wire N__27114;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27090;
    wire N__27077;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27065;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27053;
    wire N__27052;
    wire N__27051;
    wire N__27050;
    wire N__27049;
    wire N__27044;
    wire N__27043;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27023;
    wire N__27018;
    wire N__27015;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26981;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26888;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26878;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26857;
    wire N__26856;
    wire N__26853;
    wire N__26848;
    wire N__26843;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26789;
    wire N__26786;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26753;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26729;
    wire N__26728;
    wire N__26727;
    wire N__26726;
    wire N__26725;
    wire N__26722;
    wire N__26721;
    wire N__26720;
    wire N__26717;
    wire N__26716;
    wire N__26713;
    wire N__26712;
    wire N__26711;
    wire N__26702;
    wire N__26699;
    wire N__26698;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26660;
    wire N__26655;
    wire N__26654;
    wire N__26653;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26612;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26597;
    wire N__26596;
    wire N__26595;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26587;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26556;
    wire N__26553;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26535;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26524;
    wire N__26521;
    wire N__26520;
    wire N__26519;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26504;
    wire N__26497;
    wire N__26486;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26471;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26426;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26414;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26389;
    wire N__26388;
    wire N__26387;
    wire N__26386;
    wire N__26385;
    wire N__26384;
    wire N__26383;
    wire N__26382;
    wire N__26381;
    wire N__26380;
    wire N__26363;
    wire N__26362;
    wire N__26361;
    wire N__26360;
    wire N__26359;
    wire N__26358;
    wire N__26357;
    wire N__26356;
    wire N__26355;
    wire N__26354;
    wire N__26353;
    wire N__26352;
    wire N__26351;
    wire N__26350;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26342;
    wire N__26341;
    wire N__26340;
    wire N__26339;
    wire N__26338;
    wire N__26337;
    wire N__26336;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26315;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26291;
    wire N__26274;
    wire N__26271;
    wire N__26270;
    wire N__26269;
    wire N__26268;
    wire N__26267;
    wire N__26266;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26256;
    wire N__26253;
    wire N__26248;
    wire N__26245;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26221;
    wire N__26218;
    wire N__26211;
    wire N__26208;
    wire N__26203;
    wire N__26198;
    wire N__26189;
    wire N__26188;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26144;
    wire N__26143;
    wire N__26138;
    wire N__26137;
    wire N__26136;
    wire N__26135;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26120;
    wire N__26119;
    wire N__26118;
    wire N__26115;
    wire N__26114;
    wire N__26113;
    wire N__26112;
    wire N__26107;
    wire N__26106;
    wire N__26103;
    wire N__26102;
    wire N__26101;
    wire N__26100;
    wire N__26097;
    wire N__26092;
    wire N__26089;
    wire N__26088;
    wire N__26087;
    wire N__26086;
    wire N__26077;
    wire N__26076;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26055;
    wire N__26050;
    wire N__26049;
    wire N__26048;
    wire N__26045;
    wire N__26038;
    wire N__26035;
    wire N__26030;
    wire N__26027;
    wire N__26026;
    wire N__26021;
    wire N__26012;
    wire N__26007;
    wire N__26000;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25979;
    wire N__25970;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25955;
    wire N__25952;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25940;
    wire N__25939;
    wire N__25938;
    wire N__25937;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25933;
    wire N__25932;
    wire N__25929;
    wire N__25920;
    wire N__25911;
    wire N__25908;
    wire N__25903;
    wire N__25898;
    wire N__25895;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25867;
    wire N__25864;
    wire N__25861;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25743;
    wire N__25740;
    wire N__25739;
    wire N__25736;
    wire N__25727;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25673;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25640;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25609;
    wire N__25608;
    wire N__25605;
    wire N__25600;
    wire N__25599;
    wire N__25594;
    wire N__25593;
    wire N__25590;
    wire N__25589;
    wire N__25588;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25571;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25547;
    wire N__25544;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25532;
    wire N__25529;
    wire N__25528;
    wire N__25527;
    wire N__25524;
    wire N__25519;
    wire N__25514;
    wire N__25513;
    wire N__25512;
    wire N__25511;
    wire N__25508;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25490;
    wire N__25489;
    wire N__25488;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25459;
    wire N__25456;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25441;
    wire N__25438;
    wire N__25433;
    wire N__25430;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25414;
    wire N__25403;
    wire N__25400;
    wire N__25399;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25384;
    wire N__25379;
    wire N__25376;
    wire N__25375;
    wire N__25370;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25364;
    wire N__25363;
    wire N__25362;
    wire N__25361;
    wire N__25358;
    wire N__25349;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25331;
    wire N__25328;
    wire N__25327;
    wire N__25326;
    wire N__25325;
    wire N__25324;
    wire N__25323;
    wire N__25322;
    wire N__25321;
    wire N__25320;
    wire N__25317;
    wire N__25316;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25294;
    wire N__25293;
    wire N__25290;
    wire N__25273;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25228;
    wire N__25227;
    wire N__25226;
    wire N__25225;
    wire N__25222;
    wire N__25213;
    wire N__25208;
    wire N__25205;
    wire N__25204;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25186;
    wire N__25185;
    wire N__25184;
    wire N__25183;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25165;
    wire N__25154;
    wire N__25153;
    wire N__25148;
    wire N__25145;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25137;
    wire N__25134;
    wire N__25129;
    wire N__25124;
    wire N__25121;
    wire N__25120;
    wire N__25119;
    wire N__25116;
    wire N__25111;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25055;
    wire N__25054;
    wire N__25051;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25036;
    wire N__25031;
    wire N__25028;
    wire N__25027;
    wire N__25024;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24938;
    wire N__24937;
    wire N__24932;
    wire N__24929;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24914;
    wire N__24913;
    wire N__24912;
    wire N__24909;
    wire N__24904;
    wire N__24899;
    wire N__24896;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24888;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24872;
    wire N__24871;
    wire N__24868;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24853;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24802;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24749;
    wire N__24748;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24711;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24685;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24670;
    wire N__24669;
    wire N__24668;
    wire N__24665;
    wire N__24664;
    wire N__24663;
    wire N__24662;
    wire N__24659;
    wire N__24654;
    wire N__24651;
    wire N__24644;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24573;
    wire N__24570;
    wire N__24565;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24488;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24391;
    wire N__24390;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24371;
    wire N__24368;
    wire N__24367;
    wire N__24366;
    wire N__24363;
    wire N__24358;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24309;
    wire N__24306;
    wire N__24301;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24269;
    wire N__24266;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24251;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24239;
    wire N__24236;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24200;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24178;
    wire N__24177;
    wire N__24176;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24168;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24153;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24138;
    wire N__24135;
    wire N__24130;
    wire N__24119;
    wire N__24118;
    wire N__24117;
    wire N__24112;
    wire N__24109;
    wire N__24106;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24062;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24050;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24035;
    wire N__24034;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__23999;
    wire N__23998;
    wire N__23997;
    wire N__23994;
    wire N__23993;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23978;
    wire N__23975;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23960;
    wire N__23957;
    wire N__23952;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23921;
    wire N__23920;
    wire N__23919;
    wire N__23918;
    wire N__23917;
    wire N__23916;
    wire N__23913;
    wire N__23912;
    wire N__23911;
    wire N__23904;
    wire N__23901;
    wire N__23892;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23867;
    wire N__23864;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23852;
    wire N__23849;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23837;
    wire N__23834;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23822;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23792;
    wire N__23789;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23777;
    wire N__23774;
    wire N__23773;
    wire N__23772;
    wire N__23771;
    wire N__23770;
    wire N__23769;
    wire N__23766;
    wire N__23765;
    wire N__23762;
    wire N__23761;
    wire N__23758;
    wire N__23757;
    wire N__23754;
    wire N__23753;
    wire N__23752;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23730;
    wire N__23729;
    wire N__23726;
    wire N__23725;
    wire N__23722;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23710;
    wire N__23697;
    wire N__23694;
    wire N__23687;
    wire N__23684;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23669;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23642;
    wire N__23641;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23618;
    wire N__23615;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23603;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23591;
    wire N__23588;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23555;
    wire N__23552;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23531;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23516;
    wire N__23513;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23495;
    wire N__23492;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23462;
    wire N__23459;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23447;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23363;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23333;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23303;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23276;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23261;
    wire N__23258;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23239;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23204;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23189;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23165;
    wire N__23162;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23150;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23126;
    wire N__23123;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23111;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23039;
    wire N__23038;
    wire N__23037;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23026;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22970;
    wire N__22965;
    wire N__22952;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22931;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22895;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22850;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22832;
    wire N__22829;
    wire N__22828;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22808;
    wire N__22807;
    wire N__22806;
    wire N__22805;
    wire N__22804;
    wire N__22803;
    wire N__22802;
    wire N__22801;
    wire N__22796;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22780;
    wire N__22775;
    wire N__22766;
    wire N__22765;
    wire N__22764;
    wire N__22763;
    wire N__22754;
    wire N__22753;
    wire N__22752;
    wire N__22751;
    wire N__22750;
    wire N__22747;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22711;
    wire N__22708;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22693;
    wire N__22690;
    wire N__22685;
    wire N__22682;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22601;
    wire N__22600;
    wire N__22599;
    wire N__22598;
    wire N__22597;
    wire N__22596;
    wire N__22589;
    wire N__22584;
    wire N__22583;
    wire N__22580;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22559;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22548;
    wire N__22543;
    wire N__22540;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22364;
    wire N__22361;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22349;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22318;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22295;
    wire N__22292;
    wire N__22291;
    wire N__22286;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22278;
    wire N__22277;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22261;
    wire N__22260;
    wire N__22257;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22239;
    wire N__22236;
    wire N__22231;
    wire N__22226;
    wire N__22225;
    wire N__22220;
    wire N__22219;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22172;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22147;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22124;
    wire N__22123;
    wire N__22122;
    wire N__22119;
    wire N__22114;
    wire N__22109;
    wire N__22108;
    wire N__22103;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22088;
    wire N__22087;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22075;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22061;
    wire N__22058;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22027;
    wire N__22026;
    wire N__22025;
    wire N__22024;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21971;
    wire N__21964;
    wire N__21959;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21953;
    wire N__21952;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21932;
    wire N__21931;
    wire N__21926;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21911;
    wire N__21910;
    wire N__21905;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21890;
    wire N__21889;
    wire N__21888;
    wire N__21887;
    wire N__21886;
    wire N__21885;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21866;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21842;
    wire N__21837;
    wire N__21830;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21818;
    wire N__21817;
    wire N__21816;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21800;
    wire N__21797;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21755;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21743;
    wire N__21742;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21734;
    wire N__21733;
    wire N__21732;
    wire N__21731;
    wire N__21730;
    wire N__21729;
    wire N__21716;
    wire N__21713;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21683;
    wire N__21682;
    wire N__21681;
    wire N__21678;
    wire N__21677;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21669;
    wire N__21668;
    wire N__21667;
    wire N__21666;
    wire N__21665;
    wire N__21664;
    wire N__21663;
    wire N__21662;
    wire N__21659;
    wire N__21658;
    wire N__21657;
    wire N__21656;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21638;
    wire N__21633;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21611;
    wire N__21610;
    wire N__21607;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21587;
    wire N__21584;
    wire N__21575;
    wire N__21570;
    wire N__21565;
    wire N__21562;
    wire N__21551;
    wire N__21548;
    wire N__21547;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21518;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21506;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21473;
    wire N__21472;
    wire N__21467;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21452;
    wire N__21449;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21437;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21425;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21404;
    wire N__21401;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21347;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21335;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21320;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21308;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21287;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21275;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21263;
    wire N__21260;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21144;
    wire N__21139;
    wire N__21136;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21110;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21010;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20996;
    wire N__20995;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20981;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20909;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20897;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20882;
    wire N__20879;
    wire N__20878;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20864;
    wire N__20863;
    wire N__20862;
    wire N__20859;
    wire N__20854;
    wire N__20849;
    wire N__20846;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20834;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20819;
    wire N__20818;
    wire N__20817;
    wire N__20814;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20798;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20790;
    wire N__20787;
    wire N__20782;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20764;
    wire N__20763;
    wire N__20762;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20743;
    wire N__20738;
    wire N__20737;
    wire N__20736;
    wire N__20733;
    wire N__20728;
    wire N__20723;
    wire N__20722;
    wire N__20721;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20705;
    wire N__20702;
    wire N__20701;
    wire N__20700;
    wire N__20699;
    wire N__20696;
    wire N__20695;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20654;
    wire N__20651;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20633;
    wire N__20630;
    wire N__20629;
    wire N__20628;
    wire N__20625;
    wire N__20620;
    wire N__20615;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20603;
    wire N__20602;
    wire N__20599;
    wire N__20598;
    wire N__20597;
    wire N__20594;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20580;
    wire N__20577;
    wire N__20576;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20554;
    wire N__20551;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20535;
    wire N__20532;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20483;
    wire N__20482;
    wire N__20481;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20465;
    wire N__20462;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20447;
    wire N__20446;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20428;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20413;
    wire N__20412;
    wire N__20411;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20395;
    wire N__20390;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20378;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20366;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20336;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20324;
    wire N__20321;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20288;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20273;
    wire N__20270;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20251;
    wire N__20248;
    wire N__20245;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20212;
    wire N__20211;
    wire N__20210;
    wire N__20209;
    wire N__20206;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20186;
    wire N__20185;
    wire N__20184;
    wire N__20183;
    wire N__20182;
    wire N__20181;
    wire N__20178;
    wire N__20177;
    wire N__20176;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20162;
    wire N__20159;
    wire N__20154;
    wire N__20151;
    wire N__20144;
    wire N__20135;
    wire N__20134;
    wire N__20133;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20123;
    wire N__20116;
    wire N__20115;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20099;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20065;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20015;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19979;
    wire N__19976;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19928;
    wire N__19925;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19871;
    wire N__19868;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19856;
    wire N__19853;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19841;
    wire N__19838;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19756;
    wire N__19753;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19745;
    wire N__19742;
    wire N__19741;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19729;
    wire N__19726;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19706;
    wire N__19705;
    wire N__19704;
    wire N__19701;
    wire N__19700;
    wire N__19695;
    wire N__19692;
    wire N__19691;
    wire N__19690;
    wire N__19689;
    wire N__19688;
    wire N__19687;
    wire N__19686;
    wire N__19685;
    wire N__19684;
    wire N__19683;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19668;
    wire N__19667;
    wire N__19666;
    wire N__19665;
    wire N__19664;
    wire N__19649;
    wire N__19646;
    wire N__19641;
    wire N__19636;
    wire N__19627;
    wire N__19624;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19612;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19565;
    wire N__19564;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19540;
    wire N__19539;
    wire N__19536;
    wire N__19531;
    wire N__19526;
    wire N__19523;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19415;
    wire N__19414;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19400;
    wire N__19397;
    wire N__19392;
    wire N__19391;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19364;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19325;
    wire N__19320;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19259;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19241;
    wire N__19236;
    wire N__19235;
    wire N__19232;
    wire N__19227;
    wire N__19224;
    wire N__19217;
    wire N__19214;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19186;
    wire N__19183;
    wire N__19182;
    wire N__19179;
    wire N__19178;
    wire N__19177;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19151;
    wire N__19148;
    wire N__19139;
    wire N__19136;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19110;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19099;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18969;
    wire N__18964;
    wire N__18963;
    wire N__18962;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18799;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18740;
    wire N__18737;
    wire N__18736;
    wire N__18735;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18677;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18658;
    wire N__18657;
    wire N__18654;
    wire N__18649;
    wire N__18644;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18629;
    wire N__18628;
    wire N__18627;
    wire N__18624;
    wire N__18619;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18597;
    wire N__18594;
    wire N__18589;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18557;
    wire N__18554;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18539;
    wire N__18536;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18528;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18516;
    wire N__18511;
    wire N__18506;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18488;
    wire N__18485;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18471;
    wire N__18470;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18454;
    wire N__18451;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18415;
    wire N__18414;
    wire N__18413;
    wire N__18412;
    wire N__18409;
    wire N__18408;
    wire N__18405;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18389;
    wire N__18380;
    wire N__18377;
    wire N__18376;
    wire N__18375;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18364;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18348;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18338;
    wire N__18333;
    wire N__18328;
    wire N__18323;
    wire N__18320;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18316;
    wire N__18311;
    wire N__18310;
    wire N__18309;
    wire N__18308;
    wire N__18307;
    wire N__18304;
    wire N__18303;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18295;
    wire N__18294;
    wire N__18293;
    wire N__18290;
    wire N__18289;
    wire N__18282;
    wire N__18279;
    wire N__18274;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18239;
    wire N__18238;
    wire N__18237;
    wire N__18230;
    wire N__18229;
    wire N__18228;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18222;
    wire N__18211;
    wire N__18208;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18200;
    wire N__18199;
    wire N__18198;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18190;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18179;
    wire N__18178;
    wire N__18177;
    wire N__18174;
    wire N__18173;
    wire N__18166;
    wire N__18163;
    wire N__18148;
    wire N__18143;
    wire N__18140;
    wire N__18131;
    wire N__18130;
    wire N__18129;
    wire N__18128;
    wire N__18127;
    wire N__18126;
    wire N__18125;
    wire N__18124;
    wire N__18123;
    wire N__18122;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18098;
    wire N__18095;
    wire N__18090;
    wire N__18083;
    wire N__18082;
    wire N__18081;
    wire N__18080;
    wire N__18079;
    wire N__18076;
    wire N__18075;
    wire N__18074;
    wire N__18073;
    wire N__18070;
    wire N__18069;
    wire N__18066;
    wire N__18061;
    wire N__18060;
    wire N__18059;
    wire N__18058;
    wire N__18057;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18029;
    wire N__18024;
    wire N__18017;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18009;
    wire N__18008;
    wire N__18007;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17991;
    wire N__17984;
    wire N__17983;
    wire N__17982;
    wire N__17977;
    wire N__17976;
    wire N__17975;
    wire N__17972;
    wire N__17971;
    wire N__17968;
    wire N__17967;
    wire N__17966;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17954;
    wire N__17951;
    wire N__17950;
    wire N__17947;
    wire N__17946;
    wire N__17943;
    wire N__17942;
    wire N__17939;
    wire N__17938;
    wire N__17937;
    wire N__17936;
    wire N__17935;
    wire N__17932;
    wire N__17925;
    wire N__17922;
    wire N__17911;
    wire N__17904;
    wire N__17901;
    wire N__17896;
    wire N__17885;
    wire N__17884;
    wire N__17883;
    wire N__17882;
    wire N__17881;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17863;
    wire N__17862;
    wire N__17861;
    wire N__17860;
    wire N__17859;
    wire N__17858;
    wire N__17857;
    wire N__17856;
    wire N__17847;
    wire N__17846;
    wire N__17843;
    wire N__17842;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17824;
    wire N__17821;
    wire N__17812;
    wire N__17801;
    wire N__17798;
    wire N__17797;
    wire N__17796;
    wire N__17795;
    wire N__17794;
    wire N__17793;
    wire N__17788;
    wire N__17779;
    wire N__17774;
    wire N__17773;
    wire N__17772;
    wire N__17771;
    wire N__17770;
    wire N__17769;
    wire N__17768;
    wire N__17763;
    wire N__17752;
    wire N__17747;
    wire N__17746;
    wire N__17745;
    wire N__17744;
    wire N__17741;
    wire N__17740;
    wire N__17735;
    wire N__17728;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17695;
    wire N__17694;
    wire N__17693;
    wire N__17692;
    wire N__17687;
    wire N__17680;
    wire N__17677;
    wire N__17676;
    wire N__17675;
    wire N__17674;
    wire N__17673;
    wire N__17668;
    wire N__17665;
    wire N__17664;
    wire N__17663;
    wire N__17662;
    wire N__17661;
    wire N__17658;
    wire N__17657;
    wire N__17656;
    wire N__17655;
    wire N__17654;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17633;
    wire N__17630;
    wire N__17619;
    wire N__17606;
    wire N__17605;
    wire N__17604;
    wire N__17603;
    wire N__17602;
    wire N__17599;
    wire N__17592;
    wire N__17589;
    wire N__17584;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17533;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17521;
    wire N__17520;
    wire N__17515;
    wire N__17512;
    wire N__17507;
    wire N__17504;
    wire N__17503;
    wire N__17498;
    wire N__17495;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17487;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17464;
    wire N__17459;
    wire N__17458;
    wire N__17457;
    wire N__17456;
    wire N__17449;
    wire N__17446;
    wire N__17441;
    wire N__17440;
    wire N__17439;
    wire N__17436;
    wire N__17435;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17421;
    wire N__17414;
    wire N__17413;
    wire N__17412;
    wire N__17409;
    wire N__17404;
    wire N__17399;
    wire N__17396;
    wire N__17395;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17350;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17233;
    wire N__17230;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17177;
    wire N__17176;
    wire N__17173;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17158;
    wire N__17155;
    wire N__17154;
    wire N__17153;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17139;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17116;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17102;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17081;
    wire N__17078;
    wire N__17069;
    wire N__17066;
    wire N__17065;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17057;
    wire N__17056;
    wire N__17053;
    wire N__17052;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17030;
    wire N__17025;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16815;
    wire N__16814;
    wire N__16813;
    wire N__16808;
    wire N__16805;
    wire N__16804;
    wire N__16803;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16795;
    wire N__16794;
    wire N__16793;
    wire N__16792;
    wire N__16791;
    wire N__16790;
    wire N__16789;
    wire N__16784;
    wire N__16783;
    wire N__16780;
    wire N__16779;
    wire N__16778;
    wire N__16773;
    wire N__16770;
    wire N__16767;
    wire N__16752;
    wire N__16749;
    wire N__16740;
    wire N__16737;
    wire N__16732;
    wire N__16721;
    wire N__16718;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16707;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16695;
    wire N__16688;
    wire N__16687;
    wire N__16686;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16634;
    wire N__16631;
    wire N__16630;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16616;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16592;
    wire N__16583;
    wire N__16580;
    wire N__16579;
    wire N__16576;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16568;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16544;
    wire N__16535;
    wire N__16532;
    wire N__16531;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16517;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16494;
    wire N__16487;
    wire N__16484;
    wire N__16483;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16469;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16446;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16348;
    wire N__16347;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16343;
    wire N__16342;
    wire N__16341;
    wire N__16340;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16316;
    wire N__16313;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16297;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16207;
    wire N__16206;
    wire N__16199;
    wire N__16198;
    wire N__16197;
    wire N__16196;
    wire N__16193;
    wire N__16192;
    wire N__16191;
    wire N__16188;
    wire N__16187;
    wire N__16182;
    wire N__16179;
    wire N__16178;
    wire N__16177;
    wire N__16174;
    wire N__16173;
    wire N__16170;
    wire N__16165;
    wire N__16160;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16136;
    wire N__16133;
    wire N__16132;
    wire N__16131;
    wire N__16130;
    wire N__16129;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16121;
    wire N__16112;
    wire N__16109;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16091;
    wire N__16088;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16069;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16039;
    wire N__16036;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16015;
    wire N__16014;
    wire N__16013;
    wire N__16012;
    wire N__16007;
    wire N__16000;
    wire N__15999;
    wire N__15998;
    wire N__15997;
    wire N__15992;
    wire N__15991;
    wire N__15990;
    wire N__15989;
    wire N__15988;
    wire N__15987;
    wire N__15986;
    wire N__15985;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15981;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15967;
    wire N__15952;
    wire N__15951;
    wire N__15948;
    wire N__15939;
    wire N__15936;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15864;
    wire N__15861;
    wire N__15856;
    wire N__15851;
    wire N__15848;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15840;
    wire N__15837;
    wire N__15832;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15817;
    wire N__15816;
    wire N__15813;
    wire N__15808;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15719;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15656;
    wire N__15655;
    wire N__15652;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15635;
    wire N__15634;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15613;
    wire N__15608;
    wire N__15607;
    wire N__15606;
    wire N__15605;
    wire N__15604;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15572;
    wire N__15571;
    wire N__15570;
    wire N__15563;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15551;
    wire N__15550;
    wire N__15549;
    wire N__15546;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15523;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15510;
    wire N__15509;
    wire N__15508;
    wire N__15507;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15489;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15412;
    wire N__15411;
    wire N__15410;
    wire N__15401;
    wire N__15398;
    wire N__15397;
    wire N__15396;
    wire N__15395;
    wire N__15392;
    wire N__15391;
    wire N__15388;
    wire N__15379;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15337;
    wire N__15336;
    wire N__15333;
    wire N__15332;
    wire N__15323;
    wire N__15320;
    wire N__15319;
    wire N__15316;
    wire N__15315;
    wire N__15308;
    wire N__15305;
    wire N__15304;
    wire N__15301;
    wire N__15296;
    wire N__15293;
    wire N__15292;
    wire N__15291;
    wire N__15290;
    wire N__15289;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15188;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15152;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15140;
    wire N__15137;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15125;
    wire N__15122;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14992;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14971;
    wire N__14968;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14938;
    wire N__14935;
    wire N__14934;
    wire N__14931;
    wire N__14930;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14915;
    wire N__14912;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14868;
    wire N__14865;
    wire N__14864;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14843;
    wire N__14840;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14759;
    wire N__14758;
    wire N__14755;
    wire N__14754;
    wire N__14753;
    wire N__14752;
    wire N__14751;
    wire N__14750;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14738;
    wire N__14729;
    wire N__14724;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14662;
    wire N__14661;
    wire N__14658;
    wire N__14657;
    wire N__14656;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14617;
    wire N__14616;
    wire N__14615;
    wire N__14612;
    wire N__14611;
    wire N__14608;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14572;
    wire N__14571;
    wire N__14568;
    wire N__14567;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14546;
    wire N__14543;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14509;
    wire N__14504;
    wire N__14501;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14486;
    wire N__14483;
    wire N__14482;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14422;
    wire N__14419;
    wire N__14418;
    wire N__14417;
    wire N__14416;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14412;
    wire N__14405;
    wire N__14400;
    wire N__14391;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14363;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14303;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14261;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14249;
    wire N__14248;
    wire N__14243;
    wire N__14240;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14228;
    wire N__14225;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14179;
    wire N__14178;
    wire N__14177;
    wire N__14176;
    wire N__14175;
    wire N__14174;
    wire N__14173;
    wire N__14166;
    wire N__14161;
    wire N__14154;
    wire N__14147;
    wire N__14146;
    wire N__14145;
    wire N__14144;
    wire N__14143;
    wire N__14142;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14126;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14089;
    wire N__14088;
    wire N__14083;
    wire N__14080;
    wire N__14075;
    wire N__14072;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14060;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13960;
    wire N__13959;
    wire N__13958;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13946;
    wire N__13943;
    wire N__13938;
    wire N__13931;
    wire N__13930;
    wire N__13925;
    wire N__13922;
    wire N__13921;
    wire N__13916;
    wire N__13913;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13754;
    wire N__13751;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13667;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13655;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13637;
    wire N__13636;
    wire N__13633;
    wire N__13630;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13531;
    wire N__13530;
    wire N__13525;
    wire N__13522;
    wire N__13517;
    wire N__13514;
    wire N__13513;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13498;
    wire N__13497;
    wire N__13496;
    wire N__13495;
    wire N__13484;
    wire N__13481;
    wire N__13480;
    wire N__13479;
    wire N__13476;
    wire N__13475;
    wire N__13472;
    wire N__13465;
    wire N__13462;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13415;
    wire N__13412;
    wire N__13411;
    wire N__13410;
    wire N__13409;
    wire N__13408;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13392;
    wire N__13389;
    wire N__13382;
    wire N__13379;
    wire N__13378;
    wire N__13373;
    wire N__13370;
    wire N__13369;
    wire N__13366;
    wire N__13365;
    wire N__13362;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13333;
    wire N__13332;
    wire N__13331;
    wire N__13330;
    wire N__13327;
    wire N__13320;
    wire N__13317;
    wire N__13312;
    wire N__13307;
    wire N__13306;
    wire N__13305;
    wire N__13304;
    wire N__13295;
    wire N__13292;
    wire N__13291;
    wire N__13288;
    wire N__13285;
    wire N__13282;
    wire N__13277;
    wire N__13274;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13264;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13249;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire VCCG0;
    wire \Inst_eia232.Inst_transmitter.txBuffer_6 ;
    wire \Inst_eia232.Inst_transmitter.txBuffer_5 ;
    wire \Inst_eia232.Inst_transmitter.txBuffer_4 ;
    wire \Inst_eia232.Inst_transmitter.txBuffer_3 ;
    wire \Inst_eia232.Inst_transmitter.txBuffer_2 ;
    wire \Inst_eia232.Inst_transmitter.txBuffer_7 ;
    wire \Inst_eia232.Inst_transmitter.txBuffer_8 ;
    wire n234_cascade_;
    wire \Inst_eia232.Inst_transmitter.txBuffer_9 ;
    wire n234;
    wire byteDone;
    wire n9_cascade_;
    wire \Inst_eia232.Inst_transmitter.bits_3 ;
    wire \Inst_eia232.Inst_transmitter.bits_2 ;
    wire n3493;
    wire n3493_cascade_;
    wire n6749;
    wire \Inst_eia232.Inst_transmitter.bits_0 ;
    wire \Inst_eia232.Inst_transmitter.bits_1 ;
    wire n4082;
    wire \Inst_eia232.Inst_transmitter.counter_3 ;
    wire \Inst_eia232.Inst_transmitter.n2201_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.counter_4 ;
    wire \Inst_eia232.Inst_transmitter.n8642 ;
    wire \Inst_eia232.Inst_transmitter.counter_1 ;
    wire \Inst_eia232.Inst_transmitter.counter_2 ;
    wire \Inst_eia232.Inst_transmitter.n3594 ;
    wire \Inst_eia232.Inst_transmitter.n3594_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.n4719 ;
    wire n3615;
    wire \Inst_eia232.Inst_transmitter.counter_0 ;
    wire outputdata_0;
    wire outputdata_4;
    wire outputdata_5;
    wire \Inst_eia232.Inst_transmitter.txBuffer_1 ;
    wire tx_c;
    wire bfn_1_11_0_;
    wire \GENERIC_FIFO_1.n7836 ;
    wire \GENERIC_FIFO_1.n7837 ;
    wire \GENERIC_FIFO_1.n7838 ;
    wire \GENERIC_FIFO_1.n7839 ;
    wire \GENERIC_FIFO_1.n7840 ;
    wire \GENERIC_FIFO_1.n7841 ;
    wire \GENERIC_FIFO_1.n7842 ;
    wire \GENERIC_FIFO_1.n7843 ;
    wire bfn_1_12_0_;
    wire \GENERIC_FIFO_1.n7844 ;
    wire bfn_1_13_0_;
    wire \GENERIC_FIFO_1.n7827 ;
    wire \GENERIC_FIFO_1.n7828 ;
    wire \GENERIC_FIFO_1.n7829 ;
    wire \GENERIC_FIFO_1.n7830 ;
    wire \GENERIC_FIFO_1.n7831 ;
    wire \GENERIC_FIFO_1.n7832 ;
    wire \GENERIC_FIFO_1.n7833 ;
    wire \GENERIC_FIFO_1.n7834 ;
    wire bfn_1_14_0_;
    wire \GENERIC_FIFO_1.n7835 ;
    wire \GENERIC_FIFO_1.level_9_N_876_7 ;
    wire \GENERIC_FIFO_1.level_9_N_876_1 ;
    wire \GENERIC_FIFO_1.level_9_N_876_4 ;
    wire \GENERIC_FIFO_1.level_9_N_876_3 ;
    wire \GENERIC_FIFO_1.n12 ;
    wire bfn_1_15_0_;
    wire \GENERIC_FIFO_1.n11 ;
    wire \GENERIC_FIFO_1.n7818 ;
    wire \GENERIC_FIFO_1.n10 ;
    wire \GENERIC_FIFO_1.n7819 ;
    wire \GENERIC_FIFO_1.n9 ;
    wire \GENERIC_FIFO_1.n7820 ;
    wire \GENERIC_FIFO_1.n8 ;
    wire \GENERIC_FIFO_1.n7821 ;
    wire \GENERIC_FIFO_1.n7 ;
    wire \GENERIC_FIFO_1.n7822 ;
    wire \GENERIC_FIFO_1.n6 ;
    wire \GENERIC_FIFO_1.n7823 ;
    wire \GENERIC_FIFO_1.n5 ;
    wire \GENERIC_FIFO_1.n7824 ;
    wire \GENERIC_FIFO_1.n7825 ;
    wire \GENERIC_FIFO_1.n4 ;
    wire bfn_1_16_0_;
    wire \GENERIC_FIFO_1.n7826 ;
    wire \GENERIC_FIFO_1.n3 ;
    wire n4005_cascade_;
    wire dataBuffer_22;
    wire dataBuffer_30;
    wire dataBuffer_24;
    wire \Inst_eia232.Inst_transmitter.byte_0 ;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_8 ;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_0 ;
    wire \Inst_eia232.Inst_transmitter.n3571 ;
    wire dataBuffer_19;
    wire \Inst_eia232.Inst_transmitter.n8854_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.byte_3 ;
    wire dataBuffer_14;
    wire \Inst_eia232.Inst_transmitter.n1323 ;
    wire \Inst_eia232.Inst_transmitter.n3632_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.byte_6 ;
    wire dataBuffer_18;
    wire \Inst_eia232.Inst_transmitter.n8851_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.byte_2 ;
    wire \Inst_eia232.Inst_transmitter.byte_1 ;
    wire n4248_cascade_;
    wire n1336_cascade_;
    wire dataBuffer_25;
    wire \Inst_eia232.Inst_transmitter.n8847 ;
    wire n4248;
    wire n1320;
    wire n1320_cascade_;
    wire dataBuffer_28;
    wire \Inst_eia232.Inst_transmitter.n8756_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_4 ;
    wire \Inst_eia232.Inst_transmitter.byte_4 ;
    wire state_1_N_371_1_cascade_;
    wire \Inst_eia232.Inst_transmitter.n1 ;
    wire bytes_1;
    wire bytes_2;
    wire \Inst_eia232.Inst_transmitter.n9218_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.n3 ;
    wire disabled;
    wire \Inst_eia232.Inst_transmitter.n6745 ;
    wire state_1_N_371_1;
    wire \Inst_eia232.Inst_transmitter.n3652 ;
    wire bytes_0;
    wire \Inst_eia232.Inst_transmitter.n3652_cascade_ ;
    wire n1336;
    wire outputdata_1;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_1 ;
    wire outputdata_2;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_2 ;
    wire outputdata_3;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_3 ;
    wire outputdata_6;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_6 ;
    wire \Inst_eia232.Inst_transmitter.disabledBuffer_1 ;
    wire disabledGroupsReg_1;
    wire \Inst_eia232.Inst_transmitter.disabledBuffer_3 ;
    wire disabledGroupsReg_3;
    wire \Inst_eia232.Inst_transmitter.disabledBuffer_2 ;
    wire disabledGroupsReg_2;
    wire \Inst_eia232.Inst_transmitter.byte_7 ;
    wire outputdata_7;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_7 ;
    wire bfn_2_8_0_;
    wire \GENERIC_FIFO_1.n7929 ;
    wire \GENERIC_FIFO_1.n7930 ;
    wire \GENERIC_FIFO_1.n7931 ;
    wire \GENERIC_FIFO_1.n7932 ;
    wire \GENERIC_FIFO_1.n7933 ;
    wire \GENERIC_FIFO_1.n7934 ;
    wire \GENERIC_FIFO_1.n7935 ;
    wire \GENERIC_FIFO_1.n7936 ;
    wire bfn_2_9_0_;
    wire \GENERIC_FIFO_1.n7937 ;
    wire maskRegister_5;
    wire \Inst_eia232.Inst_transmitter.n6703 ;
    wire \Inst_eia232.Inst_transmitter.dataBuffer_5 ;
    wire \Inst_eia232.Inst_transmitter.byte_5 ;
    wire \GENERIC_FIFO_1.n8677_cascade_ ;
    wire \GENERIC_FIFO_1.n1396_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4743 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_0 ;
    wire \GENERIC_FIFO_1.write_pointer_8 ;
    wire \GENERIC_FIFO_1.write_pointer_9 ;
    wire \GENERIC_FIFO_1.write_pointer_7 ;
    wire \GENERIC_FIFO_1.n18_cascade_ ;
    wire \GENERIC_FIFO_1.fifo_memory_N_983 ;
    wire \GENERIC_FIFO_1.write_pointer_4 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_4 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_5 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n11 ;
    wire \GENERIC_FIFO_1.write_pointer_5 ;
    wire \GENERIC_FIFO_1.n16_cascade_ ;
    wire \GENERIC_FIFO_1.n20_adj_1274 ;
    wire \GENERIC_FIFO_1.n4721 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105 ;
    wire \GENERIC_FIFO_1.level_9_N_925_0 ;
    wire \GENERIC_FIFO_1.n24 ;
    wire bfn_2_13_0_;
    wire \GENERIC_FIFO_1.n23 ;
    wire \GENERIC_FIFO_1.n7809 ;
    wire \GENERIC_FIFO_1.n22 ;
    wire \GENERIC_FIFO_1.n7810 ;
    wire \GENERIC_FIFO_1.n21 ;
    wire \GENERIC_FIFO_1.n7811 ;
    wire \GENERIC_FIFO_1.n20 ;
    wire \GENERIC_FIFO_1.n7812 ;
    wire \GENERIC_FIFO_1.n19 ;
    wire \GENERIC_FIFO_1.n7813 ;
    wire \GENERIC_FIFO_1.n18_adj_1275 ;
    wire \GENERIC_FIFO_1.n7814 ;
    wire \GENERIC_FIFO_1.n17 ;
    wire \GENERIC_FIFO_1.n7815 ;
    wire \GENERIC_FIFO_1.n7816 ;
    wire \GENERIC_FIFO_1.n16_adj_1273 ;
    wire bfn_2_14_0_;
    wire \GENERIC_FIFO_1.n7817 ;
    wire \GENERIC_FIFO_1.n15 ;
    wire \GENERIC_FIFO_1.n8650 ;
    wire \GENERIC_FIFO_1.n8681 ;
    wire \GENERIC_FIFO_1.n78 ;
    wire \GENERIC_FIFO_1.level_9__N_900 ;
    wire \GENERIC_FIFO_1.n8654 ;
    wire \GENERIC_FIFO_1.n1418 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_6 ;
    wire \GENERIC_FIFO_1.level_9_N_876_2 ;
    wire \GENERIC_FIFO_1.level_9_N_876_6 ;
    wire \GENERIC_FIFO_1.level_9_N_876_0 ;
    wire \GENERIC_FIFO_1.level_9_N_876_8 ;
    wire \GENERIC_FIFO_1.level_9_N_876_5 ;
    wire \GENERIC_FIFO_1.n16_adj_1276_cascade_ ;
    wire \GENERIC_FIFO_1.level_9_N_876_9 ;
    wire \GENERIC_FIFO_1.n17_adj_1278 ;
    wire \GENERIC_FIFO_1.n1396 ;
    wire \GENERIC_FIFO_1.n18_adj_1277 ;
    wire \GENERIC_FIFO_1.n141_cascade_ ;
    wire \GENERIC_FIFO_1.n69 ;
    wire \Inst_eia232.Inst_receiver.n2143_cascade_ ;
    wire \Inst_eia232.Inst_receiver.bitcount_1 ;
    wire \Inst_eia232.Inst_receiver.bitcount_2 ;
    wire \Inst_eia232.Inst_receiver.bitcount_3 ;
    wire \Inst_eia232.Inst_receiver.bitcount_0 ;
    wire \Inst_eia232.Inst_receiver.n7_adj_1264_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n8769_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n6736_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n8772 ;
    wire \Inst_eia232.Inst_receiver.bytecount_2 ;
    wire \Inst_eia232.Inst_receiver.bytecount_1 ;
    wire \Inst_eia232.Inst_receiver.n8582_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n8831_cascade_ ;
    wire \Inst_eia232.Inst_transmitter.n3552 ;
    wire \Inst_eia232.xon ;
    wire \Inst_eia232.Inst_receiver.n75_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n5597 ;
    wire \Inst_eia232.Inst_receiver.n5597_cascade_ ;
    wire \Inst_eia232.xoff ;
    wire \Inst_eia232.Inst_receiver.n90_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n5498 ;
    wire cmd_6;
    wire n5698_cascade_;
    wire nstate_2_N_241_0;
    wire \Inst_eia232.Inst_receiver.n14_adj_1265 ;
    wire \Inst_eia232.Inst_receiver.n112 ;
    wire \Inst_eia232.Inst_receiver.n112_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n90 ;
    wire \GENERIC_FIFO_1.n8779 ;
    wire valueRegister_0;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n9114_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_0 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n9108 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6 ;
    wire \GENERIC_FIFO_1.n71 ;
    wire \GENERIC_FIFO_1.n70 ;
    wire \Inst_eia232.Inst_receiver.n4628 ;
    wire \Inst_eia232.Inst_transmitter.paused ;
    wire \Inst_eia232.Inst_transmitter.n4634 ;
    wire state_0;
    wire \Inst_eia232.Inst_transmitter.n2580 ;
    wire \Inst_eia232.Inst_transmitter.n8527 ;
    wire \Inst_eia232.id ;
    wire \Inst_eia232.Inst_transmitter.n971 ;
    wire state_1;
    wire \Inst_eia232.Inst_transmitter.n4712 ;
    wire \GENERIC_FIFO_1.n77 ;
    wire \GENERIC_FIFO_1.n76 ;
    wire \GENERIC_FIFO_1.n75 ;
    wire \GENERIC_FIFO_1.n74 ;
    wire \GENERIC_FIFO_1.n73 ;
    wire \GENERIC_FIFO_1.n1420 ;
    wire \GENERIC_FIFO_1.n72 ;
    wire \GENERIC_FIFO_1.n16_adj_1279_cascade_ ;
    wire \GENERIC_FIFO_1.n142 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_7 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_7 ;
    wire \GENERIC_FIFO_1.n17_adj_1280 ;
    wire \GENERIC_FIFO_1.n1421 ;
    wire \GENERIC_FIFO_1.n1423 ;
    wire writeByte;
    wire n9;
    wire \Inst_eia232.Inst_transmitter.n3608 ;
    wire \GENERIC_FIFO_1.write_pointer_0 ;
    wire \GENERIC_FIFO_1.write_pointer_1 ;
    wire \GENERIC_FIFO_1.write_pointer_2 ;
    wire \GENERIC_FIFO_1.write_pointer_3 ;
    wire \GENERIC_FIFO_1.write_pointer_6 ;
    wire \GENERIC_FIFO_1.read_pointer_0 ;
    wire \GENERIC_FIFO_1.n2 ;
    wire bfn_4_15_0_;
    wire \GENERIC_FIFO_1.n1379 ;
    wire \GENERIC_FIFO_1.n7938 ;
    wire \GENERIC_FIFO_1.n1391 ;
    wire \GENERIC_FIFO_1.n1378 ;
    wire \GENERIC_FIFO_1.n8634 ;
    wire \GENERIC_FIFO_1.n7939 ;
    wire \GENERIC_FIFO_1.n1377 ;
    wire \GENERIC_FIFO_1.n7940 ;
    wire \GENERIC_FIFO_1.n1390 ;
    wire \GENERIC_FIFO_1.n1376 ;
    wire \GENERIC_FIFO_1.n8628 ;
    wire \GENERIC_FIFO_1.n7941 ;
    wire \GENERIC_FIFO_1.n1375 ;
    wire \GENERIC_FIFO_1.n7942 ;
    wire \GENERIC_FIFO_1.n1386 ;
    wire \GENERIC_FIFO_1.n1374 ;
    wire \GENERIC_FIFO_1.n8632 ;
    wire \GENERIC_FIFO_1.n7943 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \GENERIC_FIFO_1.n7944 ;
    wire \GENERIC_FIFO_1.n7944_THRU_CRY_0_THRU_CO ;
    wire \GENERIC_FIFO_1.n1388 ;
    wire \GENERIC_FIFO_1.n1373 ;
    wire \GENERIC_FIFO_1.n8630 ;
    wire bfn_4_16_0_;
    wire \GENERIC_FIFO_1.n1372 ;
    wire \GENERIC_FIFO_1.n7945 ;
    wire \GENERIC_FIFO_1.n1383 ;
    wire \GENERIC_FIFO_1.n1371 ;
    wire \GENERIC_FIFO_1.n8638 ;
    wire \GENERIC_FIFO_1.n7946 ;
    wire \GENERIC_FIFO_1.n1392 ;
    wire \GENERIC_FIFO_1.n1392_THRU_CO ;
    wire \GENERIC_FIFO_1.n8821 ;
    wire \GENERIC_FIFO_1.read_pointer_9 ;
    wire \GENERIC_FIFO_1.n1416 ;
    wire \Inst_eia232.Inst_receiver.n8755_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n9123_cascade_ ;
    wire executePrev;
    wire \Inst_eia232.Inst_receiver.n8784 ;
    wire \Inst_eia232.Inst_receiver.n6_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n8_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n5504 ;
    wire \Inst_eia232.Inst_receiver.n8782_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n6_adj_1267 ;
    wire \Inst_eia232.Inst_receiver.n3_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n5505 ;
    wire \Inst_eia232.Inst_receiver.n3504_cascade_ ;
    wire \Inst_eia232.Inst_receiver.n3676 ;
    wire \Inst_eia232.Inst_receiver.n4767 ;
    wire \Inst_eia232.Inst_receiver.n3504 ;
    wire \Inst_eia232.Inst_receiver.n5 ;
    wire \Inst_eia232.Inst_receiver.n75 ;
    wire \Inst_eia232.Inst_receiver.n14 ;
    wire n1917;
    wire \Inst_eia232.Inst_receiver.counter_4 ;
    wire \Inst_eia232.Inst_receiver.counter_3 ;
    wire \Inst_eia232.Inst_receiver.n7_cascade_ ;
    wire \Inst_eia232.Inst_receiver.counter_1 ;
    wire \Inst_eia232.Inst_receiver.counter_0 ;
    wire \Inst_eia232.Inst_receiver.counter_2 ;
    wire \Inst_eia232.Inst_receiver.n7777 ;
    wire \Inst_eia232.Inst_receiver.n3202 ;
    wire \Inst_eia232.Inst_receiver.n1_adj_1266 ;
    wire \Inst_eia232.state_0 ;
    wire \Inst_eia232.Inst_receiver.nstate_2_N_133_1 ;
    wire \Inst_eia232.Inst_receiver.n8826 ;
    wire \Inst_eia232.Inst_prescaler.counter_4__N_38 ;
    wire \Inst_eia232.Inst_receiver.cmd_4 ;
    wire \Inst_eia232.Inst_receiver.cmd_5 ;
    wire n12;
    wire \Inst_eia232.Inst_receiver.cmd_1 ;
    wire \Inst_eia232.Inst_receiver.n3718 ;
    wire \Inst_eia232.Inst_receiver.cmd_2 ;
    wire \Inst_eia232.Inst_receiver.cmd_0 ;
    wire \Inst_eia232.Inst_receiver.cmd_3 ;
    wire \Inst_eia232.Inst_receiver.n69 ;
    wire \Inst_eia232.state_1 ;
    wire \Inst_eia232.state_2 ;
    wire \Inst_eia232.Inst_prescaler.counter_1 ;
    wire \Inst_eia232.Inst_prescaler.counter_0 ;
    wire trxClock;
    wire nstate_2__N_139_c_1;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n9096_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_cascade_ ;
    wire configRegister_23_adj_1379;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n9102_cascade_ ;
    wire valueRegister_3;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_3 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n9084_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_cascade_ ;
    wire configRegister_23_adj_1339;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n9090_cascade_ ;
    wire \Inst_core.Inst_sync.Inst_filter.n4730 ;
    wire valueRegister_2;
    wire valueRegister_5;
    wire configRegister_24;
    wire maskRegister_0_adj_1288;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4642 ;
    wire \Inst_core.Inst_sync.Inst_filter.input360_1 ;
    wire \Inst_core.Inst_sync.Inst_filter.input360_2 ;
    wire valueRegister_6;
    wire maskRegister_2;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4740 ;
    wire maskRegister_3;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4741 ;
    wire maskRegister_4;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4742 ;
    wire maskRegister_6;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4744 ;
    wire maskRegister_7;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4745 ;
    wire valueRegister_4;
    wire \GENERIC_FIFO_1.n1422 ;
    wire valueRegister_7;
    wire \Inst_core.Inst_sync.Inst_filter.n4729 ;
    wire \Inst_core.Inst_sync.Inst_filter.input360_4 ;
    wire \GENERIC_FIFO_1.n8815 ;
    wire \GENERIC_FIFO_1.read_pointer_3 ;
    wire \Inst_core.Inst_sync.Inst_filter.n4731 ;
    wire \GENERIC_FIFO_1.n1424 ;
    wire \GENERIC_FIFO_1.n1419 ;
    wire \GENERIC_FIFO_1.n8813 ;
    wire \GENERIC_FIFO_1.read_pointer_1 ;
    wire \GENERIC_FIFO_1.n8814 ;
    wire \GENERIC_FIFO_1.read_pointer_2 ;
    wire \GENERIC_FIFO_1.n1417 ;
    wire \GENERIC_FIFO_1.n8816 ;
    wire \GENERIC_FIFO_1.read_pointer_4 ;
    wire \GENERIC_FIFO_1.n8817 ;
    wire \GENERIC_FIFO_1.read_pointer_5 ;
    wire \GENERIC_FIFO_1.n8818 ;
    wire \GENERIC_FIFO_1.read_pointer_6 ;
    wire \GENERIC_FIFO_1.n8819 ;
    wire \GENERIC_FIFO_1.read_pointer_7 ;
    wire \GENERIC_FIFO_1.n141 ;
    wire \GENERIC_FIFO_1.n8820 ;
    wire \GENERIC_FIFO_1.read_pointer_8 ;
    wire \Inst_core.Inst_sync.Inst_filter.input360_0 ;
    wire \Inst_core.Inst_sync.Inst_filter.n4732 ;
    wire \Inst_core.Inst_sync.Inst_filter.input180Delay_4 ;
    wire testcnt_c_0;
    wire bfn_6_1_0_;
    wire testcnt_c_1;
    wire n7862;
    wire testcnt_c_2;
    wire n7863;
    wire testcnt_c_3;
    wire n7864;
    wire testcnt_c_4;
    wire n7865;
    wire testcnt_c_5;
    wire n7866;
    wire testcnt_c_6;
    wire n7867;
    wire n7868;
    wire testcnt_c_7;
    wire bfn_6_3_0_;
    wire configRegister_1_adj_1399;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7914 ;
    wire configRegister_2_adj_1398;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7915 ;
    wire configRegister_3_adj_1397;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7916 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7917 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7918 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7919 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7920 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7921 ;
    wire configRegister_8_adj_1392;
    wire bfn_6_4_0_;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7922 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7923 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7924 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7925 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7926 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7927 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7928 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15 ;
    wire \Inst_eia232.Inst_receiver.n7_adj_1264 ;
    wire \Inst_eia232.Inst_receiver.n957 ;
    wire \Inst_eia232.Inst_receiver.bytecount_0 ;
    wire \Inst_eia232.Inst_receiver.n3557 ;
    wire \Inst_eia232.Inst_receiver.n8376 ;
    wire maskRegister_6_adj_1362;
    wire maskRegister_7_adj_1361;
    wire maskRegister_4_adj_1364;
    wire configRegister_6_adj_1394;
    wire maskRegister_3_adj_1365;
    wire configRegister_7_adj_1393;
    wire valueRegister_0_adj_1296;
    wire \Inst_core.Inst_sync.Inst_filter.input360_3 ;
    wire configRegister_0_adj_1400;
    wire configRegister_20_adj_1342;
    wire configRegister_4_adj_1396;
    wire cmd_39;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4641 ;
    wire configRegister_21_adj_1381;
    wire wrtrigval_0;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1 ;
    wire valueRegister_1;
    wire configRegister_26;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_1 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n9078 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_cascade_ ;
    wire configRegister_21_adj_1301;
    wire configRegister_23_adj_1299;
    wire configRegister_22_adj_1300;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n9072_cascade_ ;
    wire configRegister_20_adj_1302;
    wire configRegister_24_adj_1298;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0 ;
    wire maskRegister_1_adj_1287;
    wire maskRegister_2_adj_1286;
    wire maskRegister_3_adj_1285;
    wire maskRegister_5_adj_1283;
    wire \Inst_core.Inst_sync.filteredInput_2 ;
    wire \Inst_core.Inst_sync.n2789_cascade_ ;
    wire syncedInput_2;
    wire \Inst_core.Inst_sync.demuxedInput_6 ;
    wire \Inst_core.Inst_sync.filteredInput_6 ;
    wire maskRegister_4_adj_1284;
    wire \Inst_core.Inst_sync.Inst_filter.n4637 ;
    wire maskRegister_1;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4739 ;
    wire \Inst_core.Inst_sync.Inst_filter.input180Delay_7 ;
    wire \Inst_core.Inst_sync.filteredInput_5 ;
    wire \Inst_core.Inst_sync.n9063_cascade_ ;
    wire syncedInput_5;
    wire \Inst_core.Inst_sync.synchronizedInput_4 ;
    wire \Inst_core.Inst_sync.filteredInput_4 ;
    wire \Inst_core.Inst_sync.demuxedInput_4 ;
    wire \Inst_core.Inst_sync.n9057_cascade_ ;
    wire syncedInput_4;
    wire \Inst_core.Inst_sync.Inst_filter.input180Delay_6 ;
    wire \Inst_core.Inst_sync.Inst_filter.n4734 ;
    wire \Inst_core.Inst_sync.Inst_filter.input180Delay_5 ;
    wire \Inst_core.Inst_sync.Inst_filter.n4733 ;
    wire input_c_4;
    wire \Inst_core.Inst_sync.synchronizedInput180_4 ;
    wire \INVInst_core.Inst_sync.synchronizedInput180_i4C_net ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4765 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n25_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n27 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n26 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4766 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n28 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n28 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n25_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n27 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n26 ;
    wire valueRegister_6_adj_1370;
    wire configRegister_5_adj_1395;
    wire valueRegister_7_adj_1369;
    wire configRegister_11_adj_1389;
    wire configRegister_10_adj_1390;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_7 ;
    wire configRegister_15_adj_1385;
    wire configRegister_24_adj_1378;
    wire \Inst_eia232.Inst_transmitter.n4246 ;
    wire n4005;
    wire disabledGroupsReg_0;
    wire \Inst_eia232.Inst_transmitter.disabledBuffer_0 ;
    wire configRegister_22_adj_1380;
    wire configRegister_23;
    wire wrtrigmask_0;
    wire maskRegister_0;
    wire configRegister_20_adj_1382;
    wire configRegister_22_adj_1340;
    wire configRegister_21;
    wire wrtrigmask_1;
    wire configRegister_21_adj_1341;
    wire wrFlags;
    wire cmd_32;
    wire configRegister_20;
    wire valueRegister_1_adj_1295;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_1 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4746 ;
    wire fwd_15;
    wire \Inst_core.Inst_controller.n22_cascade_ ;
    wire fwd_6;
    wire \Inst_core.Inst_controller.n4_adj_986_cascade_ ;
    wire fwd_5;
    wire \Inst_core.Inst_controller.n4_adj_987_cascade_ ;
    wire \Inst_core.Inst_controller.n8486 ;
    wire \Inst_core.Inst_sync.demuxedInput_0 ;
    wire syncedInput_3;
    wire syncedInput_7;
    wire valueRegister_7_adj_1329;
    wire \Inst_core.Inst_sync.filteredInput_1 ;
    wire \Inst_core.Inst_sync.filteredInput_3 ;
    wire \Inst_core.Inst_sync.n2791 ;
    wire \Inst_core.Inst_sync.filteredInput_0 ;
    wire \Inst_core.Inst_sync.n2793 ;
    wire flagInverted;
    wire flagFilter;
    wire \Inst_core.Inst_sync.demuxedInput_1 ;
    wire \Inst_core.Inst_sync.n2787 ;
    wire \Inst_core.Inst_sync.Inst_filter.input360_5 ;
    wire syncedInput_6;
    wire \Inst_core.Inst_sync.Inst_filter.input360_6 ;
    wire \Inst_core.Inst_sync.demuxedInput_7 ;
    wire \Inst_core.Inst_sync.demuxedInput_2 ;
    wire \Inst_core.Inst_sync.demuxedInput_5 ;
    wire \Inst_core.Inst_sync.n9117 ;
    wire \Inst_core.Inst_sync.demuxedInput_3 ;
    wire \Inst_core.Inst_sync.synchronizedInput_5 ;
    wire \Inst_core.Inst_sync.n2566 ;
    wire \Inst_core.Inst_sync.n2564 ;
    wire \Inst_core.Inst_sync.n9129 ;
    wire \Inst_core.Inst_sync.synchronizedInput_6 ;
    wire input_c_0;
    wire \Inst_core.Inst_sync.synchronizedInput180_0 ;
    wire input_c_1;
    wire \Inst_core.Inst_sync.synchronizedInput180_1 ;
    wire input_c_2;
    wire \Inst_core.Inst_sync.synchronizedInput180_2 ;
    wire input_c_3;
    wire \Inst_core.Inst_sync.synchronizedInput180_3 ;
    wire input_c_6;
    wire \Inst_core.Inst_sync.synchronizedInput180_6 ;
    wire input_c_5;
    wire \Inst_core.Inst_sync.synchronizedInput180_5 ;
    wire \Inst_core.Inst_sync.synchronizedInput180_7 ;
    wire \INVInst_core.Inst_sync.synchronizedInput180_i0C_net ;
    wire \Inst_core.n8518_cascade_ ;
    wire valueRegister_7_adj_1289;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_7 ;
    wire memoryOut_7;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n8808_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n3 ;
    wire \Inst_core.n1639_cascade_ ;
    wire \Inst_core.n9054 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0 ;
    wire bfn_8_2_0_;
    wire configRegister_1_adj_1359;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7899 ;
    wire configRegister_2_adj_1358;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7900 ;
    wire configRegister_3_adj_1357;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7901 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7902 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7903 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7904 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7905 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7906 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8 ;
    wire bfn_8_3_0_;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7907 ;
    wire configRegister_10_adj_1350;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7908 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7909 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7910 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7911 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7912 ;
    wire \Inst_core.n1639 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7913 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4114 ;
    wire \Inst_core.configRegister_27 ;
    wire configRegister_7_adj_1353;
    wire configRegister_11_adj_1349;
    wire configRegister_12_adj_1388;
    wire configRegister_5_adj_1355;
    wire configRegister_14_adj_1346;
    wire configRegister_9_adj_1351;
    wire configRegister_8_adj_1352;
    wire cmd_16;
    wire configRegister_15_adj_1345;
    wire wrtrigmask_3;
    wire configRegister_9_adj_1391;
    wire cmd_38;
    wire \Inst_core.Inst_controller.fwd_14 ;
    wire cmd_30;
    wire configRegister_22;
    wire cmd_33;
    wire cmd_37;
    wire cmd_36;
    wire configRegister_6_adj_1354;
    wire valueRegister_5_adj_1291;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4750 ;
    wire bwd_11;
    wire bwd_8;
    wire fwd_11;
    wire fwd_4;
    wire \Inst_core.Inst_controller.n18_cascade_ ;
    wire \Inst_core.Inst_controller.n21 ;
    wire fwd_13;
    wire fwd_9;
    wire \Inst_core.Inst_controller.n15 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4 ;
    wire valueRegister_4_adj_1292;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4749 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_5 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_7 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_4 ;
    wire fwd_12;
    wire fwd_1;
    wire \Inst_core.Inst_controller.n13 ;
    wire bwd_10;
    wire \Inst_core.Inst_controller.n14 ;
    wire fwd_8;
    wire \Inst_core.Inst_controller.n11 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n14 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n11 ;
    wire cmd_29;
    wire syncedInput_0;
    wire syncedInput_1;
    wire valueRegister_4_adj_1332;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4756 ;
    wire \Inst_core.Inst_sampler.n31_adj_995_cascade_ ;
    wire divider_9;
    wire divider_7;
    wire \Inst_core.Inst_sampler.n29 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_7 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_4 ;
    wire valueRegister_5_adj_1331;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_5 ;
    wire divider_15;
    wire divider_13;
    wire divider_16;
    wire \Inst_core.Inst_sampler.n32 ;
    wire divider_14;
    wire \Inst_core.Inst_sampler.n8596_cascade_ ;
    wire \Inst_core.Inst_sampler.n8590 ;
    wire valueRegister_1_adj_1335;
    wire divider_20;
    wire divider_21;
    wire \Inst_core.Inst_sampler.n8598 ;
    wire \Inst_core.Inst_sampler.n8602 ;
    wire \Inst_core.Inst_sampler.n8600_cascade_ ;
    wire \Inst_core.Inst_sampler.n8604 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelL16 ;
    wire configRegister_24_adj_1338;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_7 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n8844_cascade_ ;
    wire \Inst_core.Inst_decoder.n6 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n9052 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n1765 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n667 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n667_cascade_ ;
    wire \Inst_core.n31_adj_1174 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n100_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n656 ;
    wire \Inst_core.n8518 ;
    wire \Inst_core.state_1_adj_1134 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n657 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n554 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n22_cascade_ ;
    wire \Inst_core.n8515_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n451 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n760 ;
    wire \Inst_core.n31 ;
    wire cmd_18;
    wire configRegister_13_adj_1347;
    wire configRegister_14_adj_1386;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5 ;
    wire memoryOut_5;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n2_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n100 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n553 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n100_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n2_cascade_ ;
    wire configRegister_17_adj_1383;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n100 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n100_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n759 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n770 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.state_1 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n770_cascade_ ;
    wire \Inst_core.n6713 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4076 ;
    wire configRegister_17_adj_1303;
    wire configRegister_4_adj_1356;
    wire maskRegister_5_adj_1363;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4764 ;
    wire configRegister_12_adj_1348;
    wire \Inst_core.arm ;
    wire maskRegister_5_adj_1323;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4757 ;
    wire maskRegister_6_adj_1322;
    wire maskRegister_7_adj_1321;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4759 ;
    wire maskRegister_0_adj_1368;
    wire maskRegister_1_adj_1367;
    wire maskRegister_2_adj_1366;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7_adj_996 ;
    wire flagDemux;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register ;
    wire valueRegister_5_adj_1371;
    wire configRegister_13_adj_1387;
    wire wrtrigcfg_3;
    wire configRegister_16_adj_1384;
    wire configRegister_16_adj_1304;
    wire cmd_17;
    wire cmd_28;
    wire fwd_3;
    wire bwd_9;
    wire \Inst_core.Inst_controller.n24 ;
    wire \Inst_core.Inst_controller.n22_adj_988_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3 ;
    wire valueRegister_3_adj_1293;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_3 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4748 ;
    wire bwd_6;
    wire bwd_5;
    wire \Inst_core.Inst_controller.n23 ;
    wire bwd_3;
    wire bwd_4;
    wire \Inst_core.Inst_controller.n21_adj_989 ;
    wire cmd_11;
    wire cmd_15;
    wire bwd_7;
    wire fwd_10;
    wire wrtrigmask_2;
    wire maskRegister_4_adj_1324;
    wire \Inst_core.Inst_sync.filteredInput_7 ;
    wire \Inst_core.Inst_sync.Inst_filter.n4735 ;
    wire maskRegister_7_adj_1281;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4752 ;
    wire maskRegister_0_adj_1328;
    wire maskRegister_1_adj_1327;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4753 ;
    wire maskRegister_2_adj_1326;
    wire maskRegister_3_adj_1325;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6 ;
    wire valueRegister_6_adj_1330;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_6 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4758 ;
    wire divider_4;
    wire \Inst_core.Inst_sampler.n30 ;
    wire \Inst_core.Inst_sampler.n8592 ;
    wire divider_2;
    wire divider_10;
    wire divider_8;
    wire divider_17;
    wire \Inst_core.Inst_sampler.n8588 ;
    wire bfn_9_14_0_;
    wire \Inst_core.Inst_sampler.n7948 ;
    wire \Inst_core.Inst_sampler.n7949 ;
    wire \Inst_core.Inst_sampler.n7950 ;
    wire \Inst_core.Inst_sampler.counter_4 ;
    wire \Inst_core.Inst_sampler.n7951 ;
    wire \Inst_core.Inst_sampler.n7952 ;
    wire \Inst_core.Inst_sampler.n7953 ;
    wire \Inst_core.Inst_sampler.counter_7 ;
    wire \Inst_core.Inst_sampler.n7954 ;
    wire \Inst_core.Inst_sampler.n7955 ;
    wire \Inst_core.Inst_sampler.counter_8 ;
    wire bfn_9_15_0_;
    wire \Inst_core.Inst_sampler.counter_9 ;
    wire \Inst_core.Inst_sampler.n7956 ;
    wire \Inst_core.Inst_sampler.counter_10 ;
    wire \Inst_core.Inst_sampler.n7957 ;
    wire \Inst_core.Inst_sampler.n7958 ;
    wire \Inst_core.Inst_sampler.n7959 ;
    wire \Inst_core.Inst_sampler.counter_13 ;
    wire \Inst_core.Inst_sampler.n7960 ;
    wire \Inst_core.Inst_sampler.counter_14 ;
    wire \Inst_core.Inst_sampler.n7961 ;
    wire \Inst_core.Inst_sampler.counter_15 ;
    wire \Inst_core.Inst_sampler.n7962 ;
    wire \Inst_core.Inst_sampler.n7963 ;
    wire \Inst_core.Inst_sampler.counter_16 ;
    wire bfn_9_16_0_;
    wire \Inst_core.Inst_sampler.counter_17 ;
    wire \Inst_core.Inst_sampler.n7964 ;
    wire \Inst_core.Inst_sampler.n7965 ;
    wire \Inst_core.Inst_sampler.counter_19 ;
    wire \Inst_core.Inst_sampler.n7966 ;
    wire \Inst_core.Inst_sampler.counter_20 ;
    wire \Inst_core.Inst_sampler.n7967 ;
    wire \Inst_core.Inst_sampler.counter_21 ;
    wire \Inst_core.Inst_sampler.n7968 ;
    wire \Inst_core.Inst_sampler.n7969 ;
    wire \Inst_core.Inst_sampler.n7970 ;
    wire \Inst_core.Inst_sampler.n1700 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n8622 ;
    wire cmd_35;
    wire configRegister_0_adj_1360;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4 ;
    wire memoryOut_4;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4763 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_5 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_7 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_6 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_4 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n11 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n6675_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n564 ;
    wire \Inst_core.n8837 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.state_1 ;
    wire configRegister_0_adj_1320;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n9055 ;
    wire bfn_11_4_0_;
    wire configRegister_1_adj_1319;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7884 ;
    wire configRegister_2_adj_1318;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7885 ;
    wire configRegister_3_adj_1317;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7886 ;
    wire configRegister_4_adj_1316;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7887 ;
    wire configRegister_5_adj_1315;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7888 ;
    wire configRegister_6_adj_1314;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7889 ;
    wire configRegister_7_adj_1313;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7890 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7891 ;
    wire configRegister_8_adj_1312;
    wire bfn_11_5_0_;
    wire configRegister_9_adj_1311;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7892 ;
    wire configRegister_10_adj_1310;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7893 ;
    wire configRegister_11_adj_1309;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7894 ;
    wire configRegister_12_adj_1308;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7895 ;
    wire configRegister_13_adj_1307;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7896 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7897 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n1662 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n7898 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4144 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4761 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n2_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n100 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n100_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n450 ;
    wire \Inst_core.Inst_trigger.levelReg_0 ;
    wire configRegister_17_adj_1343;
    wire \Inst_core.Inst_trigger.levelReg_1 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n99 ;
    wire valueRegister_4_adj_1372;
    wire configRegister_15_adj_1305;
    wire bwd_15;
    wire configRegister_17;
    wire cmd_21;
    wire wrtrigcfg_1;
    wire configRegister_14_adj_1306;
    wire cmd_12;
    wire fwd_7;
    wire maskRegister_6_adj_1282;
    wire cmd_31;
    wire cmd_10;
    wire valueRegister_2_adj_1374;
    wire cmd_25;
    wire wrtrigval_2;
    wire cmd_22;
    wire cmd_26;
    wire cmd_27;
    wire divider_19;
    wire bwd_2;
    wire bwd_13;
    wire \Inst_core.Inst_controller.n18_adj_990 ;
    wire \Inst_core.Inst_controller.n20 ;
    wire \Inst_core.Inst_controller.n17_cascade_ ;
    wire \Inst_core.Inst_controller.n30 ;
    wire \Inst_core.Inst_controller.n29_cascade_ ;
    wire \Inst_core.Inst_controller.n6693 ;
    wire \Inst_core.Inst_controller.bwd_14 ;
    wire \Inst_core.Inst_controller.n19 ;
    wire valueRegister_2_adj_1294;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4747 ;
    wire memoryOut_6;
    wire configRegister_26_adj_1297;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_6 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n4751 ;
    wire fwd_0;
    wire fwd_2;
    wire \Inst_core.Inst_controller.n16 ;
    wire debugleds_c_1;
    wire \Inst_core.n4_cascade_ ;
    wire \Inst_core.Inst_controller.n3907_cascade_ ;
    wire memoryOut_2;
    wire valueRegister_2_adj_1334;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4754 ;
    wire divider_11;
    wire \Inst_core.Inst_sampler.counter_23 ;
    wire \Inst_core.Inst_sampler.counter_11 ;
    wire \Inst_core.Inst_sampler.counter_2 ;
    wire \Inst_core.Inst_sampler.n8606 ;
    wire \Inst_core.Inst_sampler.n3_cascade_ ;
    wire divider_23;
    wire \Inst_core.Inst_sampler.n8618 ;
    wire \Inst_core.Inst_sampler.n8656_cascade_ ;
    wire divider_1;
    wire \Inst_core.Inst_sampler.counter_18 ;
    wire divider_18;
    wire \Inst_core.Inst_sampler.counter_1 ;
    wire \Inst_core.Inst_sampler.n28 ;
    wire \Inst_core.Inst_sampler.n27_cascade_ ;
    wire divider_6;
    wire \Inst_core.Inst_sampler.counter_3 ;
    wire divider_3;
    wire \Inst_core.Inst_sampler.counter_6 ;
    wire \Inst_core.Inst_sampler.n26 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3 ;
    wire valueRegister_3_adj_1333;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4755 ;
    wire divider_0;
    wire \Inst_core.Inst_sampler.counter_12 ;
    wire divider_12;
    wire \Inst_core.Inst_sampler.counter_0 ;
    wire \Inst_core.Inst_sampler.n25 ;
    wire \Inst_core.Inst_sync.Inst_filter.input360_7 ;
    wire input_c_7;
    wire \Inst_core.Inst_sync.synchronizedInput_7 ;
    wire cmd_13;
    wire \Inst_core.Inst_sampler.n35 ;
    wire \Inst_core.Inst_sampler.n36 ;
    wire \Inst_core.Inst_sampler.n33 ;
    wire wrDivider;
    wire \Inst_core.Inst_sampler.n8669 ;
    wire \Inst_core.Inst_sampler.n8671 ;
    wire \Inst_core.Inst_sampler.n8673 ;
    wire \Inst_core.Inst_sampler.n8687 ;
    wire valueRegister_0_adj_1336;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n4643 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_1 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_3 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_0 ;
    wire \Inst_core.Inst_trigger.stages_2__Inst_stage.n7 ;
    wire divider_5;
    wire \Inst_core.Inst_sampler.counter_22 ;
    wire divider_22;
    wire \Inst_core.Inst_sampler.counter_5 ;
    wire \Inst_core.Inst_sampler.n34 ;
    wire \Inst_core.Inst_sampler.n44 ;
    wire \Inst_core.Inst_sampler.n43 ;
    wire \Inst_core.Inst_sampler.n45 ;
    wire ready50_N_581;
    wire \Inst_core.configRegister_27_adj_1196 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n8626 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4 ;
    wire memoryOut_0;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4645 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_2 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_0 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7_adj_1000 ;
    wire \Inst_core.Inst_trigger.configRegister_27 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n8521_cascade_ ;
    wire \Inst_core.n3670 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n7 ;
    wire \Inst_core.Inst_trigger.stageRun_0 ;
    wire \Inst_core.Inst_trigger.stageRun_3 ;
    wire \Inst_core.stageRun_2 ;
    wire \Inst_core.stageRun_1 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n8753_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n461 ;
    wire \Inst_core.state_1 ;
    wire valueRegister_3_adj_1373;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3 ;
    wire memoryOut_3;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_3 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4762 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n28 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n25_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n31 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n27 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8 ;
    wire \Inst_core.Inst_trigger.stages_1__Inst_stage.n26 ;
    wire configRegister_0;
    wire \Inst_core.n9053 ;
    wire bfn_12_5_0_;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7869 ;
    wire configRegister_2;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7870 ;
    wire configRegister_3;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7871 ;
    wire configRegister_4;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7872 ;
    wire configRegister_5;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7873 ;
    wire configRegister_6;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7874 ;
    wire configRegister_7;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7875 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7876 ;
    wire configRegister_8;
    wire bfn_12_6_0_;
    wire configRegister_9;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7877 ;
    wire configRegister_10;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7878 ;
    wire configRegister_11;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7879 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7880 ;
    wire configRegister_13;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7881 ;
    wire configRegister_14;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7882 ;
    wire \Inst_core.n1705 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n7883 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n4044 ;
    wire valueRegister_1_adj_1375;
    wire memoryOut_1;
    wire configRegister_26_adj_1377;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_1 ;
    wire \Inst_core.Inst_trigger.stages_3__Inst_stage.n4760 ;
    wire \Inst_core.Inst_trigger.stageMatch_2 ;
    wire \Inst_core.Inst_trigger.stageMatch_3 ;
    wire \Inst_core.Inst_trigger.stageMatch_1 ;
    wire \Inst_core.Inst_trigger.stageMatch_0 ;
    wire \Inst_core.Inst_trigger.levelReg_1__N_590 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n28 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n25_cascade_ ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n27 ;
    wire \Inst_core.n31_adj_1132 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3 ;
    wire \Inst_core.Inst_trigger.stages_0__Inst_stage.n26 ;
    wire configRegister_1;
    wire configRegister_16;
    wire n3753;
    wire n1;
    wire cmd_19;
    wire wrtrigval_1;
    wire cmd_14;
    wire valueRegister_6_adj_1290;
    wire configRegister_12;
    wire cmd_9;
    wire bwd_1;
    wire wrtrigcfg_0;
    wire cmd_23;
    wire configRegister_15;
    wire cmd_24;
    wire configRegister_16_adj_1344;
    wire wrtrigval_3;
    wire valueRegister_0_adj_1376;
    wire cmd_8;
    wire bwd_0;
    wire wrtrigcfg_2;
    wire cmd_34;
    wire configRegister_26_adj_1337;
    wire wrsize;
    wire cmd_20;
    wire bwd_12;
    wire \Inst_core.nstate_1_N_831_0 ;
    wire \Inst_core.Inst_controller.n321 ;
    wire \Inst_core.Inst_controller.nstate_1_N_827_1 ;
    wire \Inst_core.resetCmd ;
    wire debugleds_c_0;
    wire busy;
    wire \Inst_core.Inst_controller.nstate_1_N_825_0 ;
    wire \Inst_core.Inst_controller.n320 ;
    wire \Inst_core.Inst_controller.nstate_1_N_829_0 ;
    wire \Inst_core.Inst_controller.n2717 ;
    wire sampleReady;
    wire \Inst_core.n318 ;
    wire \Inst_core.Inst_controller.n2717_cascade_ ;
    wire send;
    wire \Inst_core.Inst_controller.n2 ;
    wire \Inst_core.Inst_controller.counter_0 ;
    wire bfn_12_12_0_;
    wire \Inst_core.Inst_controller.counter_1 ;
    wire \Inst_core.Inst_controller.n7845 ;
    wire \Inst_core.Inst_controller.counter_2 ;
    wire \Inst_core.Inst_controller.n7846 ;
    wire \Inst_core.Inst_controller.counter_3 ;
    wire \Inst_core.Inst_controller.n7847 ;
    wire \Inst_core.Inst_controller.counter_4 ;
    wire \Inst_core.Inst_controller.n7848 ;
    wire \Inst_core.Inst_controller.counter_5 ;
    wire \Inst_core.Inst_controller.n7849 ;
    wire \Inst_core.Inst_controller.counter_6 ;
    wire \Inst_core.Inst_controller.n7850 ;
    wire \Inst_core.Inst_controller.counter_7 ;
    wire \Inst_core.Inst_controller.n7851 ;
    wire \Inst_core.Inst_controller.n7852 ;
    wire \Inst_core.Inst_controller.counter_8 ;
    wire bfn_12_13_0_;
    wire \Inst_core.Inst_controller.counter_9 ;
    wire \Inst_core.Inst_controller.n7853 ;
    wire \Inst_core.Inst_controller.counter_10 ;
    wire \Inst_core.Inst_controller.n7854 ;
    wire \Inst_core.Inst_controller.counter_11 ;
    wire \Inst_core.Inst_controller.n7855 ;
    wire \Inst_core.Inst_controller.counter_12 ;
    wire \Inst_core.Inst_controller.n7856 ;
    wire \Inst_core.Inst_controller.counter_13 ;
    wire \Inst_core.Inst_controller.n7857 ;
    wire \Inst_core.Inst_controller.counter_14 ;
    wire \Inst_core.Inst_controller.n7858 ;
    wire \Inst_core.Inst_controller.counter_15 ;
    wire \Inst_core.Inst_controller.n7859 ;
    wire \Inst_core.Inst_controller.n7860 ;
    wire \Inst_core.Inst_controller.counter_16 ;
    wire bfn_12_14_0_;
    wire \Inst_core.Inst_controller.n7861 ;
    wire \Inst_core.Inst_controller.counter_17 ;
    wire _gnd_net_;
    wire xtalClock_c;
    wire \Inst_core.Inst_controller.n3907 ;
    wire \Inst_core.Inst_controller.n4691 ;

    defparam \GENERIC_FIFO_1.fifo_memory0_physical .WRITE_MODE=2;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .READ_MODE=2;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory0_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \GENERIC_FIFO_1.fifo_memory0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,outputdata_7,dangling_wire_2,dangling_wire_3,dangling_wire_4,outputdata_6,dangling_wire_5,dangling_wire_6,dangling_wire_7,outputdata_5,dangling_wire_8,dangling_wire_9,dangling_wire_10,outputdata_4,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__15362,N__15761,N__15782,N__16367,N__16394,N__16409,N__16424,N__16439,N__15887,N__15257}),
            .WADDR({dangling_wire_13,N__14627,N__14672,N__14579,N__17120,N__14879,N__14948,N__16487,N__16535,N__16583,N__16634}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__23046,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__30462,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__25513,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__28076,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__37486),
            .RE(N__17350),
            .WCLKE(),
            .WCLK(N__37487),
            .WE(N__14992));
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .WRITE_MODE=2;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .READ_MODE=2;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \GENERIC_FIFO_1.fifo_memory1_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \GENERIC_FIFO_1.fifo_memory1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,outputdata_3,dangling_wire_44,dangling_wire_45,dangling_wire_46,outputdata_2,dangling_wire_47,dangling_wire_48,dangling_wire_49,outputdata_1,dangling_wire_50,dangling_wire_51,dangling_wire_52,outputdata_0,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__15356,N__15755,N__15776,N__16361,N__16388,N__16403,N__16418,N__16433,N__15881,N__15251}),
            .WADDR({dangling_wire_55,N__14621,N__14666,N__14573,N__17112,N__14872,N__14942,N__16479,N__16527,N__16576,N__16626}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__32337,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__30935,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__33651,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__31817,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__37500),
            .RE(N__17354),
            .WCLKE(),
            .WCLK(N__37499),
            .WE(N__14991));
    PRE_IO_GBUF xtalClock_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__38004),
            .GLOBALBUFFEROUTPUT(xtalClock_c));
    defparam xtalClock_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam xtalClock_pad_iopad.PULLUP=1'b0;
    IO_PAD xtalClock_pad_iopad (
            .OE(N__38006),
            .DIN(N__38005),
            .DOUT(N__38004),
            .PACKAGEPIN(xtalClock));
    defparam xtalClock_pad_preio.PIN_TYPE=6'b000001;
    defparam xtalClock_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO xtalClock_pad_preio (
            .PADOEN(N__38006),
            .PADOUT(N__38005),
            .PADIN(N__38004),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam debugleds_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam debugleds_pad_0_iopad.PULLUP=1'b0;
    IO_PAD debugleds_pad_0_iopad (
            .OE(N__37995),
            .DIN(N__37994),
            .DOUT(N__37993),
            .PACKAGEPIN(debugleds[0]));
    defparam debugleds_pad_0_preio.PIN_TYPE=6'b011001;
    defparam debugleds_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO debugleds_pad_0_preio (
            .PADOEN(N__37995),
            .PADOUT(N__37994),
            .PADIN(N__37993),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36737),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam debugleds_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam debugleds_pad_1_iopad.PULLUP=1'b0;
    IO_PAD debugleds_pad_1_iopad (
            .OE(N__37986),
            .DIN(N__37985),
            .DOUT(N__37984),
            .PACKAGEPIN(debugleds[1]));
    defparam debugleds_pad_1_preio.PIN_TYPE=6'b011001;
    defparam debugleds_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO debugleds_pad_1_preio (
            .PADOEN(N__37986),
            .PADOUT(N__37985),
            .PADIN(N__37984),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30155),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_0_iopad.PULLUP=1'b0;
    IO_PAD input_pad_0_iopad (
            .OE(N__37977),
            .DIN(N__37976),
            .DOUT(N__37975),
            .PACKAGEPIN(\input [0]));
    defparam input_pad_0_preio.PIN_TYPE=6'b000001;
    defparam input_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_0_preio (
            .PADOEN(N__37977),
            .PADOUT(N__37976),
            .PADIN(N__37975),
            .CLOCKENABLE(),
            .DIN0(input_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_1_iopad.PULLUP=1'b0;
    IO_PAD input_pad_1_iopad (
            .OE(N__37968),
            .DIN(N__37967),
            .DOUT(N__37966),
            .PACKAGEPIN(\input [1]));
    defparam input_pad_1_preio.PIN_TYPE=6'b000001;
    defparam input_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_1_preio (
            .PADOEN(N__37968),
            .PADOUT(N__37967),
            .PADIN(N__37966),
            .CLOCKENABLE(),
            .DIN0(input_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_2_iopad.PULLUP=1'b0;
    IO_PAD input_pad_2_iopad (
            .OE(N__37959),
            .DIN(N__37958),
            .DOUT(N__37957),
            .PACKAGEPIN(\input [2]));
    defparam input_pad_2_preio.PIN_TYPE=6'b000001;
    defparam input_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_2_preio (
            .PADOEN(N__37959),
            .PADOUT(N__37958),
            .PADIN(N__37957),
            .CLOCKENABLE(),
            .DIN0(input_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_3_iopad.PULLUP=1'b0;
    IO_PAD input_pad_3_iopad (
            .OE(N__37950),
            .DIN(N__37949),
            .DOUT(N__37948),
            .PACKAGEPIN(\input [3]));
    defparam input_pad_3_preio.PIN_TYPE=6'b000001;
    defparam input_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_3_preio (
            .PADOEN(N__37950),
            .PADOUT(N__37949),
            .PADIN(N__37948),
            .CLOCKENABLE(),
            .DIN0(input_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_4_iopad.PULLUP=1'b0;
    IO_PAD input_pad_4_iopad (
            .OE(N__37941),
            .DIN(N__37940),
            .DOUT(N__37939),
            .PACKAGEPIN(\input [4]));
    defparam input_pad_4_preio.PIN_TYPE=6'b000001;
    defparam input_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_4_preio (
            .PADOEN(N__37941),
            .PADOUT(N__37940),
            .PADIN(N__37939),
            .CLOCKENABLE(),
            .DIN0(input_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_5_iopad.PULLUP=1'b0;
    IO_PAD input_pad_5_iopad (
            .OE(N__37932),
            .DIN(N__37931),
            .DOUT(N__37930),
            .PACKAGEPIN(\input [5]));
    defparam input_pad_5_preio.PIN_TYPE=6'b000001;
    defparam input_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_5_preio (
            .PADOEN(N__37932),
            .PADOUT(N__37931),
            .PADIN(N__37930),
            .CLOCKENABLE(),
            .DIN0(input_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_6_iopad.PULLUP=1'b0;
    IO_PAD input_pad_6_iopad (
            .OE(N__37923),
            .DIN(N__37922),
            .DOUT(N__37921),
            .PACKAGEPIN(\input [6]));
    defparam input_pad_6_preio.PIN_TYPE=6'b000001;
    defparam input_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_6_preio (
            .PADOEN(N__37923),
            .PADOUT(N__37922),
            .PADIN(N__37921),
            .CLOCKENABLE(),
            .DIN0(input_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam input_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam input_pad_7_iopad.PULLUP=1'b0;
    IO_PAD input_pad_7_iopad (
            .OE(N__37914),
            .DIN(N__37913),
            .DOUT(N__37912),
            .PACKAGEPIN(\input [7]));
    defparam input_pad_7_preio.PIN_TYPE=6'b000001;
    defparam input_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO input_pad_7_preio (
            .PADOEN(N__37914),
            .PADOUT(N__37913),
            .PADIN(N__37912),
            .CLOCKENABLE(),
            .DIN0(input_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam nstate_2__N_139_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam nstate_2__N_139_pad_1_iopad.PULLUP=1'b0;
    IO_PAD nstate_2__N_139_pad_1_iopad (
            .OE(N__37905),
            .DIN(N__37904),
            .DOUT(N__37903),
            .PACKAGEPIN(rx));
    defparam nstate_2__N_139_pad_1_preio.PIN_TYPE=6'b000001;
    defparam nstate_2__N_139_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO nstate_2__N_139_pad_1_preio (
            .PADOEN(N__37905),
            .PADOUT(N__37904),
            .PADIN(N__37903),
            .CLOCKENABLE(),
            .DIN0(nstate_2__N_139_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ready50_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ready50_pad_iopad.PULLUP=1'b0;
    IO_PAD ready50_pad_iopad (
            .OE(N__37896),
            .DIN(N__37895),
            .DOUT(N__37894),
            .PACKAGEPIN(ready50));
    defparam ready50_pad_preio.PIN_TYPE=6'b010101;
    defparam ready50_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ready50_pad_preio (
            .PADOEN(N__37896),
            .PADOUT(N__37895),
            .PADIN(N__37894),
            .CLOCKENABLE(N__32228),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31956),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__37621),
            .OUTPUTENABLE());
    defparam testcnt_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_0_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_0_iopad (
            .OE(N__37887),
            .DIN(N__37886),
            .DOUT(N__37885),
            .PACKAGEPIN(testcnt[0]));
    defparam testcnt_pad_0_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_0_preio (
            .PADOEN(N__37887),
            .PADOUT(N__37886),
            .PADIN(N__37885),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19487),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam testcnt_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_1_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_1_iopad (
            .OE(N__37878),
            .DIN(N__37877),
            .DOUT(N__37876),
            .PACKAGEPIN(testcnt[1]));
    defparam testcnt_pad_1_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_1_preio (
            .PADOEN(N__37878),
            .PADOUT(N__37877),
            .PADIN(N__37876),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19910),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam testcnt_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_2_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_2_iopad (
            .OE(N__37869),
            .DIN(N__37868),
            .DOUT(N__37867),
            .PACKAGEPIN(testcnt[2]));
    defparam testcnt_pad_2_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_2_preio (
            .PADOEN(N__37869),
            .PADOUT(N__37868),
            .PADIN(N__37867),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19889),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam testcnt_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_3_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_3_iopad (
            .OE(N__37860),
            .DIN(N__37859),
            .DOUT(N__37858),
            .PACKAGEPIN(testcnt[3]));
    defparam testcnt_pad_3_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_3_preio (
            .PADOEN(N__37860),
            .PADOUT(N__37859),
            .PADIN(N__37858),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19868),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam testcnt_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_4_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_4_iopad (
            .OE(N__37851),
            .DIN(N__37850),
            .DOUT(N__37849),
            .PACKAGEPIN(testcnt[4]));
    defparam testcnt_pad_4_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_4_preio (
            .PADOEN(N__37851),
            .PADOUT(N__37850),
            .PADIN(N__37849),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19853),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam testcnt_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_5_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_5_iopad (
            .OE(N__37842),
            .DIN(N__37841),
            .DOUT(N__37840),
            .PACKAGEPIN(testcnt[5]));
    defparam testcnt_pad_5_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_5_preio (
            .PADOEN(N__37842),
            .PADOUT(N__37841),
            .PADIN(N__37840),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19838),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam testcnt_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_6_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_6_iopad (
            .OE(N__37833),
            .DIN(N__37832),
            .DOUT(N__37831),
            .PACKAGEPIN(testcnt[6]));
    defparam testcnt_pad_6_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_6_preio (
            .PADOEN(N__37833),
            .PADOUT(N__37832),
            .PADIN(N__37831),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19823),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam testcnt_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam testcnt_pad_7_iopad.PULLUP=1'b0;
    IO_PAD testcnt_pad_7_iopad (
            .OE(N__37824),
            .DIN(N__37823),
            .DOUT(N__37822),
            .PACKAGEPIN(testcnt[7]));
    defparam testcnt_pad_7_preio.PIN_TYPE=6'b011001;
    defparam testcnt_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO testcnt_pad_7_preio (
            .PADOEN(N__37824),
            .PADOUT(N__37823),
            .PADIN(N__37822),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19799),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_pad_iopad.PULLUP=1'b0;
    IO_PAD tx_pad_iopad (
            .OE(N__37815),
            .DIN(N__37814),
            .DOUT(N__37813),
            .PACKAGEPIN(tx));
    defparam tx_pad_preio.PIN_TYPE=6'b011001;
    defparam tx_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_pad_preio (
            .PADOEN(N__37815),
            .PADOUT(N__37814),
            .PADIN(N__37813),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13559),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__9296 (
            .O(N__37796),
            .I(N__37790));
    InMux I__9295 (
            .O(N__37795),
            .I(N__37790));
    LocalMux I__9294 (
            .O(N__37790),
            .I(N__37786));
    InMux I__9293 (
            .O(N__37789),
            .I(N__37783));
    Span4Mux_h I__9292 (
            .O(N__37786),
            .I(N__37780));
    LocalMux I__9291 (
            .O(N__37783),
            .I(\Inst_core.Inst_controller.counter_12 ));
    Odrv4 I__9290 (
            .O(N__37780),
            .I(\Inst_core.Inst_controller.counter_12 ));
    InMux I__9289 (
            .O(N__37775),
            .I(\Inst_core.Inst_controller.n7856 ));
    InMux I__9288 (
            .O(N__37772),
            .I(N__37766));
    InMux I__9287 (
            .O(N__37771),
            .I(N__37766));
    LocalMux I__9286 (
            .O(N__37766),
            .I(N__37762));
    InMux I__9285 (
            .O(N__37765),
            .I(N__37759));
    Span4Mux_v I__9284 (
            .O(N__37762),
            .I(N__37756));
    LocalMux I__9283 (
            .O(N__37759),
            .I(\Inst_core.Inst_controller.counter_13 ));
    Odrv4 I__9282 (
            .O(N__37756),
            .I(\Inst_core.Inst_controller.counter_13 ));
    InMux I__9281 (
            .O(N__37751),
            .I(\Inst_core.Inst_controller.n7857 ));
    InMux I__9280 (
            .O(N__37748),
            .I(N__37742));
    InMux I__9279 (
            .O(N__37747),
            .I(N__37742));
    LocalMux I__9278 (
            .O(N__37742),
            .I(N__37738));
    InMux I__9277 (
            .O(N__37741),
            .I(N__37735));
    Span4Mux_h I__9276 (
            .O(N__37738),
            .I(N__37732));
    LocalMux I__9275 (
            .O(N__37735),
            .I(\Inst_core.Inst_controller.counter_14 ));
    Odrv4 I__9274 (
            .O(N__37732),
            .I(\Inst_core.Inst_controller.counter_14 ));
    InMux I__9273 (
            .O(N__37727),
            .I(\Inst_core.Inst_controller.n7858 ));
    InMux I__9272 (
            .O(N__37724),
            .I(N__37720));
    InMux I__9271 (
            .O(N__37723),
            .I(N__37716));
    LocalMux I__9270 (
            .O(N__37720),
            .I(N__37713));
    InMux I__9269 (
            .O(N__37719),
            .I(N__37710));
    LocalMux I__9268 (
            .O(N__37716),
            .I(N__37705));
    Span4Mux_h I__9267 (
            .O(N__37713),
            .I(N__37705));
    LocalMux I__9266 (
            .O(N__37710),
            .I(\Inst_core.Inst_controller.counter_15 ));
    Odrv4 I__9265 (
            .O(N__37705),
            .I(\Inst_core.Inst_controller.counter_15 ));
    InMux I__9264 (
            .O(N__37700),
            .I(\Inst_core.Inst_controller.n7859 ));
    InMux I__9263 (
            .O(N__37697),
            .I(N__37693));
    InMux I__9262 (
            .O(N__37696),
            .I(N__37690));
    LocalMux I__9261 (
            .O(N__37693),
            .I(N__37687));
    LocalMux I__9260 (
            .O(N__37690),
            .I(N__37681));
    Span4Mux_h I__9259 (
            .O(N__37687),
            .I(N__37681));
    InMux I__9258 (
            .O(N__37686),
            .I(N__37678));
    Span4Mux_h I__9257 (
            .O(N__37681),
            .I(N__37675));
    LocalMux I__9256 (
            .O(N__37678),
            .I(\Inst_core.Inst_controller.counter_16 ));
    Odrv4 I__9255 (
            .O(N__37675),
            .I(\Inst_core.Inst_controller.counter_16 ));
    InMux I__9254 (
            .O(N__37670),
            .I(bfn_12_14_0_));
    InMux I__9253 (
            .O(N__37667),
            .I(\Inst_core.Inst_controller.n7861 ));
    InMux I__9252 (
            .O(N__37664),
            .I(N__37660));
    InMux I__9251 (
            .O(N__37663),
            .I(N__37657));
    LocalMux I__9250 (
            .O(N__37660),
            .I(N__37653));
    LocalMux I__9249 (
            .O(N__37657),
            .I(N__37650));
    InMux I__9248 (
            .O(N__37656),
            .I(N__37647));
    Span4Mux_h I__9247 (
            .O(N__37653),
            .I(N__37644));
    Span4Mux_h I__9246 (
            .O(N__37650),
            .I(N__37641));
    LocalMux I__9245 (
            .O(N__37647),
            .I(N__37636));
    Span4Mux_v I__9244 (
            .O(N__37644),
            .I(N__37636));
    Span4Mux_h I__9243 (
            .O(N__37641),
            .I(N__37633));
    Odrv4 I__9242 (
            .O(N__37636),
            .I(\Inst_core.Inst_controller.counter_17 ));
    Odrv4 I__9241 (
            .O(N__37633),
            .I(\Inst_core.Inst_controller.counter_17 ));
    ClkMux I__9240 (
            .O(N__37628),
            .I(N__37163));
    ClkMux I__9239 (
            .O(N__37627),
            .I(N__37163));
    ClkMux I__9238 (
            .O(N__37626),
            .I(N__37163));
    ClkMux I__9237 (
            .O(N__37625),
            .I(N__37163));
    ClkMux I__9236 (
            .O(N__37624),
            .I(N__37163));
    ClkMux I__9235 (
            .O(N__37623),
            .I(N__37163));
    ClkMux I__9234 (
            .O(N__37622),
            .I(N__37163));
    ClkMux I__9233 (
            .O(N__37621),
            .I(N__37163));
    ClkMux I__9232 (
            .O(N__37620),
            .I(N__37163));
    ClkMux I__9231 (
            .O(N__37619),
            .I(N__37163));
    ClkMux I__9230 (
            .O(N__37618),
            .I(N__37163));
    ClkMux I__9229 (
            .O(N__37617),
            .I(N__37163));
    ClkMux I__9228 (
            .O(N__37616),
            .I(N__37163));
    ClkMux I__9227 (
            .O(N__37615),
            .I(N__37163));
    ClkMux I__9226 (
            .O(N__37614),
            .I(N__37163));
    ClkMux I__9225 (
            .O(N__37613),
            .I(N__37163));
    ClkMux I__9224 (
            .O(N__37612),
            .I(N__37163));
    ClkMux I__9223 (
            .O(N__37611),
            .I(N__37163));
    ClkMux I__9222 (
            .O(N__37610),
            .I(N__37163));
    ClkMux I__9221 (
            .O(N__37609),
            .I(N__37163));
    ClkMux I__9220 (
            .O(N__37608),
            .I(N__37163));
    ClkMux I__9219 (
            .O(N__37607),
            .I(N__37163));
    ClkMux I__9218 (
            .O(N__37606),
            .I(N__37163));
    ClkMux I__9217 (
            .O(N__37605),
            .I(N__37163));
    ClkMux I__9216 (
            .O(N__37604),
            .I(N__37163));
    ClkMux I__9215 (
            .O(N__37603),
            .I(N__37163));
    ClkMux I__9214 (
            .O(N__37602),
            .I(N__37163));
    ClkMux I__9213 (
            .O(N__37601),
            .I(N__37163));
    ClkMux I__9212 (
            .O(N__37600),
            .I(N__37163));
    ClkMux I__9211 (
            .O(N__37599),
            .I(N__37163));
    ClkMux I__9210 (
            .O(N__37598),
            .I(N__37163));
    ClkMux I__9209 (
            .O(N__37597),
            .I(N__37163));
    ClkMux I__9208 (
            .O(N__37596),
            .I(N__37163));
    ClkMux I__9207 (
            .O(N__37595),
            .I(N__37163));
    ClkMux I__9206 (
            .O(N__37594),
            .I(N__37163));
    ClkMux I__9205 (
            .O(N__37593),
            .I(N__37163));
    ClkMux I__9204 (
            .O(N__37592),
            .I(N__37163));
    ClkMux I__9203 (
            .O(N__37591),
            .I(N__37163));
    ClkMux I__9202 (
            .O(N__37590),
            .I(N__37163));
    ClkMux I__9201 (
            .O(N__37589),
            .I(N__37163));
    ClkMux I__9200 (
            .O(N__37588),
            .I(N__37163));
    ClkMux I__9199 (
            .O(N__37587),
            .I(N__37163));
    ClkMux I__9198 (
            .O(N__37586),
            .I(N__37163));
    ClkMux I__9197 (
            .O(N__37585),
            .I(N__37163));
    ClkMux I__9196 (
            .O(N__37584),
            .I(N__37163));
    ClkMux I__9195 (
            .O(N__37583),
            .I(N__37163));
    ClkMux I__9194 (
            .O(N__37582),
            .I(N__37163));
    ClkMux I__9193 (
            .O(N__37581),
            .I(N__37163));
    ClkMux I__9192 (
            .O(N__37580),
            .I(N__37163));
    ClkMux I__9191 (
            .O(N__37579),
            .I(N__37163));
    ClkMux I__9190 (
            .O(N__37578),
            .I(N__37163));
    ClkMux I__9189 (
            .O(N__37577),
            .I(N__37163));
    ClkMux I__9188 (
            .O(N__37576),
            .I(N__37163));
    ClkMux I__9187 (
            .O(N__37575),
            .I(N__37163));
    ClkMux I__9186 (
            .O(N__37574),
            .I(N__37163));
    ClkMux I__9185 (
            .O(N__37573),
            .I(N__37163));
    ClkMux I__9184 (
            .O(N__37572),
            .I(N__37163));
    ClkMux I__9183 (
            .O(N__37571),
            .I(N__37163));
    ClkMux I__9182 (
            .O(N__37570),
            .I(N__37163));
    ClkMux I__9181 (
            .O(N__37569),
            .I(N__37163));
    ClkMux I__9180 (
            .O(N__37568),
            .I(N__37163));
    ClkMux I__9179 (
            .O(N__37567),
            .I(N__37163));
    ClkMux I__9178 (
            .O(N__37566),
            .I(N__37163));
    ClkMux I__9177 (
            .O(N__37565),
            .I(N__37163));
    ClkMux I__9176 (
            .O(N__37564),
            .I(N__37163));
    ClkMux I__9175 (
            .O(N__37563),
            .I(N__37163));
    ClkMux I__9174 (
            .O(N__37562),
            .I(N__37163));
    ClkMux I__9173 (
            .O(N__37561),
            .I(N__37163));
    ClkMux I__9172 (
            .O(N__37560),
            .I(N__37163));
    ClkMux I__9171 (
            .O(N__37559),
            .I(N__37163));
    ClkMux I__9170 (
            .O(N__37558),
            .I(N__37163));
    ClkMux I__9169 (
            .O(N__37557),
            .I(N__37163));
    ClkMux I__9168 (
            .O(N__37556),
            .I(N__37163));
    ClkMux I__9167 (
            .O(N__37555),
            .I(N__37163));
    ClkMux I__9166 (
            .O(N__37554),
            .I(N__37163));
    ClkMux I__9165 (
            .O(N__37553),
            .I(N__37163));
    ClkMux I__9164 (
            .O(N__37552),
            .I(N__37163));
    ClkMux I__9163 (
            .O(N__37551),
            .I(N__37163));
    ClkMux I__9162 (
            .O(N__37550),
            .I(N__37163));
    ClkMux I__9161 (
            .O(N__37549),
            .I(N__37163));
    ClkMux I__9160 (
            .O(N__37548),
            .I(N__37163));
    ClkMux I__9159 (
            .O(N__37547),
            .I(N__37163));
    ClkMux I__9158 (
            .O(N__37546),
            .I(N__37163));
    ClkMux I__9157 (
            .O(N__37545),
            .I(N__37163));
    ClkMux I__9156 (
            .O(N__37544),
            .I(N__37163));
    ClkMux I__9155 (
            .O(N__37543),
            .I(N__37163));
    ClkMux I__9154 (
            .O(N__37542),
            .I(N__37163));
    ClkMux I__9153 (
            .O(N__37541),
            .I(N__37163));
    ClkMux I__9152 (
            .O(N__37540),
            .I(N__37163));
    ClkMux I__9151 (
            .O(N__37539),
            .I(N__37163));
    ClkMux I__9150 (
            .O(N__37538),
            .I(N__37163));
    ClkMux I__9149 (
            .O(N__37537),
            .I(N__37163));
    ClkMux I__9148 (
            .O(N__37536),
            .I(N__37163));
    ClkMux I__9147 (
            .O(N__37535),
            .I(N__37163));
    ClkMux I__9146 (
            .O(N__37534),
            .I(N__37163));
    ClkMux I__9145 (
            .O(N__37533),
            .I(N__37163));
    ClkMux I__9144 (
            .O(N__37532),
            .I(N__37163));
    ClkMux I__9143 (
            .O(N__37531),
            .I(N__37163));
    ClkMux I__9142 (
            .O(N__37530),
            .I(N__37163));
    ClkMux I__9141 (
            .O(N__37529),
            .I(N__37163));
    ClkMux I__9140 (
            .O(N__37528),
            .I(N__37163));
    ClkMux I__9139 (
            .O(N__37527),
            .I(N__37163));
    ClkMux I__9138 (
            .O(N__37526),
            .I(N__37163));
    ClkMux I__9137 (
            .O(N__37525),
            .I(N__37163));
    ClkMux I__9136 (
            .O(N__37524),
            .I(N__37163));
    ClkMux I__9135 (
            .O(N__37523),
            .I(N__37163));
    ClkMux I__9134 (
            .O(N__37522),
            .I(N__37163));
    ClkMux I__9133 (
            .O(N__37521),
            .I(N__37163));
    ClkMux I__9132 (
            .O(N__37520),
            .I(N__37163));
    ClkMux I__9131 (
            .O(N__37519),
            .I(N__37163));
    ClkMux I__9130 (
            .O(N__37518),
            .I(N__37163));
    ClkMux I__9129 (
            .O(N__37517),
            .I(N__37163));
    ClkMux I__9128 (
            .O(N__37516),
            .I(N__37163));
    ClkMux I__9127 (
            .O(N__37515),
            .I(N__37163));
    ClkMux I__9126 (
            .O(N__37514),
            .I(N__37163));
    ClkMux I__9125 (
            .O(N__37513),
            .I(N__37163));
    ClkMux I__9124 (
            .O(N__37512),
            .I(N__37163));
    ClkMux I__9123 (
            .O(N__37511),
            .I(N__37163));
    ClkMux I__9122 (
            .O(N__37510),
            .I(N__37163));
    ClkMux I__9121 (
            .O(N__37509),
            .I(N__37163));
    ClkMux I__9120 (
            .O(N__37508),
            .I(N__37163));
    ClkMux I__9119 (
            .O(N__37507),
            .I(N__37163));
    ClkMux I__9118 (
            .O(N__37506),
            .I(N__37163));
    ClkMux I__9117 (
            .O(N__37505),
            .I(N__37163));
    ClkMux I__9116 (
            .O(N__37504),
            .I(N__37163));
    ClkMux I__9115 (
            .O(N__37503),
            .I(N__37163));
    ClkMux I__9114 (
            .O(N__37502),
            .I(N__37163));
    ClkMux I__9113 (
            .O(N__37501),
            .I(N__37163));
    ClkMux I__9112 (
            .O(N__37500),
            .I(N__37163));
    ClkMux I__9111 (
            .O(N__37499),
            .I(N__37163));
    ClkMux I__9110 (
            .O(N__37498),
            .I(N__37163));
    ClkMux I__9109 (
            .O(N__37497),
            .I(N__37163));
    ClkMux I__9108 (
            .O(N__37496),
            .I(N__37163));
    ClkMux I__9107 (
            .O(N__37495),
            .I(N__37163));
    ClkMux I__9106 (
            .O(N__37494),
            .I(N__37163));
    ClkMux I__9105 (
            .O(N__37493),
            .I(N__37163));
    ClkMux I__9104 (
            .O(N__37492),
            .I(N__37163));
    ClkMux I__9103 (
            .O(N__37491),
            .I(N__37163));
    ClkMux I__9102 (
            .O(N__37490),
            .I(N__37163));
    ClkMux I__9101 (
            .O(N__37489),
            .I(N__37163));
    ClkMux I__9100 (
            .O(N__37488),
            .I(N__37163));
    ClkMux I__9099 (
            .O(N__37487),
            .I(N__37163));
    ClkMux I__9098 (
            .O(N__37486),
            .I(N__37163));
    ClkMux I__9097 (
            .O(N__37485),
            .I(N__37163));
    ClkMux I__9096 (
            .O(N__37484),
            .I(N__37163));
    ClkMux I__9095 (
            .O(N__37483),
            .I(N__37163));
    ClkMux I__9094 (
            .O(N__37482),
            .I(N__37163));
    ClkMux I__9093 (
            .O(N__37481),
            .I(N__37163));
    ClkMux I__9092 (
            .O(N__37480),
            .I(N__37163));
    ClkMux I__9091 (
            .O(N__37479),
            .I(N__37163));
    ClkMux I__9090 (
            .O(N__37478),
            .I(N__37163));
    ClkMux I__9089 (
            .O(N__37477),
            .I(N__37163));
    ClkMux I__9088 (
            .O(N__37476),
            .I(N__37163));
    ClkMux I__9087 (
            .O(N__37475),
            .I(N__37163));
    ClkMux I__9086 (
            .O(N__37474),
            .I(N__37163));
    GlobalMux I__9085 (
            .O(N__37163),
            .I(N__37160));
    gio2CtrlBuf I__9084 (
            .O(N__37160),
            .I(xtalClock_c));
    CEMux I__9083 (
            .O(N__37157),
            .I(N__37153));
    CEMux I__9082 (
            .O(N__37156),
            .I(N__37149));
    LocalMux I__9081 (
            .O(N__37153),
            .I(N__37146));
    CEMux I__9080 (
            .O(N__37152),
            .I(N__37143));
    LocalMux I__9079 (
            .O(N__37149),
            .I(N__37140));
    Span4Mux_s0_h I__9078 (
            .O(N__37146),
            .I(N__37135));
    LocalMux I__9077 (
            .O(N__37143),
            .I(N__37135));
    Span4Mux_v I__9076 (
            .O(N__37140),
            .I(N__37132));
    Span4Mux_v I__9075 (
            .O(N__37135),
            .I(N__37127));
    Span4Mux_s0_h I__9074 (
            .O(N__37132),
            .I(N__37127));
    Odrv4 I__9073 (
            .O(N__37127),
            .I(\Inst_core.Inst_controller.n3907 ));
    SRMux I__9072 (
            .O(N__37124),
            .I(N__37121));
    LocalMux I__9071 (
            .O(N__37121),
            .I(N__37118));
    Span4Mux_s1_h I__9070 (
            .O(N__37118),
            .I(N__37113));
    SRMux I__9069 (
            .O(N__37117),
            .I(N__37110));
    SRMux I__9068 (
            .O(N__37116),
            .I(N__37107));
    Odrv4 I__9067 (
            .O(N__37113),
            .I(\Inst_core.Inst_controller.n4691 ));
    LocalMux I__9066 (
            .O(N__37110),
            .I(\Inst_core.Inst_controller.n4691 ));
    LocalMux I__9065 (
            .O(N__37107),
            .I(\Inst_core.Inst_controller.n4691 ));
    InMux I__9064 (
            .O(N__37100),
            .I(N__37095));
    InMux I__9063 (
            .O(N__37099),
            .I(N__37092));
    InMux I__9062 (
            .O(N__37098),
            .I(N__37089));
    LocalMux I__9061 (
            .O(N__37095),
            .I(\Inst_core.Inst_controller.counter_4 ));
    LocalMux I__9060 (
            .O(N__37092),
            .I(\Inst_core.Inst_controller.counter_4 ));
    LocalMux I__9059 (
            .O(N__37089),
            .I(\Inst_core.Inst_controller.counter_4 ));
    InMux I__9058 (
            .O(N__37082),
            .I(\Inst_core.Inst_controller.n7848 ));
    InMux I__9057 (
            .O(N__37079),
            .I(N__37075));
    InMux I__9056 (
            .O(N__37078),
            .I(N__37072));
    LocalMux I__9055 (
            .O(N__37075),
            .I(N__37066));
    LocalMux I__9054 (
            .O(N__37072),
            .I(N__37066));
    InMux I__9053 (
            .O(N__37071),
            .I(N__37063));
    Span4Mux_h I__9052 (
            .O(N__37066),
            .I(N__37060));
    LocalMux I__9051 (
            .O(N__37063),
            .I(\Inst_core.Inst_controller.counter_5 ));
    Odrv4 I__9050 (
            .O(N__37060),
            .I(\Inst_core.Inst_controller.counter_5 ));
    InMux I__9049 (
            .O(N__37055),
            .I(\Inst_core.Inst_controller.n7849 ));
    InMux I__9048 (
            .O(N__37052),
            .I(N__37048));
    InMux I__9047 (
            .O(N__37051),
            .I(N__37045));
    LocalMux I__9046 (
            .O(N__37048),
            .I(N__37039));
    LocalMux I__9045 (
            .O(N__37045),
            .I(N__37039));
    InMux I__9044 (
            .O(N__37044),
            .I(N__37036));
    Span4Mux_h I__9043 (
            .O(N__37039),
            .I(N__37033));
    LocalMux I__9042 (
            .O(N__37036),
            .I(\Inst_core.Inst_controller.counter_6 ));
    Odrv4 I__9041 (
            .O(N__37033),
            .I(\Inst_core.Inst_controller.counter_6 ));
    InMux I__9040 (
            .O(N__37028),
            .I(\Inst_core.Inst_controller.n7850 ));
    InMux I__9039 (
            .O(N__37025),
            .I(N__37021));
    InMux I__9038 (
            .O(N__37024),
            .I(N__37018));
    LocalMux I__9037 (
            .O(N__37021),
            .I(N__37015));
    LocalMux I__9036 (
            .O(N__37018),
            .I(N__37011));
    Span4Mux_v I__9035 (
            .O(N__37015),
            .I(N__37008));
    InMux I__9034 (
            .O(N__37014),
            .I(N__37005));
    Span4Mux_v I__9033 (
            .O(N__37011),
            .I(N__37002));
    Span4Mux_h I__9032 (
            .O(N__37008),
            .I(N__36999));
    LocalMux I__9031 (
            .O(N__37005),
            .I(\Inst_core.Inst_controller.counter_7 ));
    Odrv4 I__9030 (
            .O(N__37002),
            .I(\Inst_core.Inst_controller.counter_7 ));
    Odrv4 I__9029 (
            .O(N__36999),
            .I(\Inst_core.Inst_controller.counter_7 ));
    InMux I__9028 (
            .O(N__36992),
            .I(\Inst_core.Inst_controller.n7851 ));
    InMux I__9027 (
            .O(N__36989),
            .I(N__36985));
    InMux I__9026 (
            .O(N__36988),
            .I(N__36982));
    LocalMux I__9025 (
            .O(N__36985),
            .I(N__36979));
    LocalMux I__9024 (
            .O(N__36982),
            .I(N__36975));
    Span4Mux_h I__9023 (
            .O(N__36979),
            .I(N__36972));
    InMux I__9022 (
            .O(N__36978),
            .I(N__36969));
    Span4Mux_h I__9021 (
            .O(N__36975),
            .I(N__36966));
    Span4Mux_h I__9020 (
            .O(N__36972),
            .I(N__36963));
    LocalMux I__9019 (
            .O(N__36969),
            .I(\Inst_core.Inst_controller.counter_8 ));
    Odrv4 I__9018 (
            .O(N__36966),
            .I(\Inst_core.Inst_controller.counter_8 ));
    Odrv4 I__9017 (
            .O(N__36963),
            .I(\Inst_core.Inst_controller.counter_8 ));
    InMux I__9016 (
            .O(N__36956),
            .I(bfn_12_13_0_));
    InMux I__9015 (
            .O(N__36953),
            .I(N__36947));
    InMux I__9014 (
            .O(N__36952),
            .I(N__36947));
    LocalMux I__9013 (
            .O(N__36947),
            .I(N__36943));
    InMux I__9012 (
            .O(N__36946),
            .I(N__36940));
    Span4Mux_h I__9011 (
            .O(N__36943),
            .I(N__36937));
    LocalMux I__9010 (
            .O(N__36940),
            .I(\Inst_core.Inst_controller.counter_9 ));
    Odrv4 I__9009 (
            .O(N__36937),
            .I(\Inst_core.Inst_controller.counter_9 ));
    InMux I__9008 (
            .O(N__36932),
            .I(\Inst_core.Inst_controller.n7853 ));
    InMux I__9007 (
            .O(N__36929),
            .I(N__36925));
    InMux I__9006 (
            .O(N__36928),
            .I(N__36922));
    LocalMux I__9005 (
            .O(N__36925),
            .I(N__36916));
    LocalMux I__9004 (
            .O(N__36922),
            .I(N__36916));
    InMux I__9003 (
            .O(N__36921),
            .I(N__36913));
    Span4Mux_v I__9002 (
            .O(N__36916),
            .I(N__36910));
    LocalMux I__9001 (
            .O(N__36913),
            .I(\Inst_core.Inst_controller.counter_10 ));
    Odrv4 I__9000 (
            .O(N__36910),
            .I(\Inst_core.Inst_controller.counter_10 ));
    InMux I__8999 (
            .O(N__36905),
            .I(\Inst_core.Inst_controller.n7854 ));
    InMux I__8998 (
            .O(N__36902),
            .I(N__36898));
    InMux I__8997 (
            .O(N__36901),
            .I(N__36895));
    LocalMux I__8996 (
            .O(N__36898),
            .I(N__36889));
    LocalMux I__8995 (
            .O(N__36895),
            .I(N__36889));
    InMux I__8994 (
            .O(N__36894),
            .I(N__36886));
    Span4Mux_h I__8993 (
            .O(N__36889),
            .I(N__36883));
    LocalMux I__8992 (
            .O(N__36886),
            .I(\Inst_core.Inst_controller.counter_11 ));
    Odrv4 I__8991 (
            .O(N__36883),
            .I(\Inst_core.Inst_controller.counter_11 ));
    InMux I__8990 (
            .O(N__36878),
            .I(\Inst_core.Inst_controller.n7855 ));
    SRMux I__8989 (
            .O(N__36875),
            .I(N__36868));
    CascadeMux I__8988 (
            .O(N__36874),
            .I(N__36861));
    CascadeMux I__8987 (
            .O(N__36873),
            .I(N__36855));
    InMux I__8986 (
            .O(N__36872),
            .I(N__36851));
    InMux I__8985 (
            .O(N__36871),
            .I(N__36848));
    LocalMux I__8984 (
            .O(N__36868),
            .I(N__36845));
    CascadeMux I__8983 (
            .O(N__36867),
            .I(N__36841));
    InMux I__8982 (
            .O(N__36866),
            .I(N__36838));
    SRMux I__8981 (
            .O(N__36865),
            .I(N__36835));
    SRMux I__8980 (
            .O(N__36864),
            .I(N__36832));
    InMux I__8979 (
            .O(N__36861),
            .I(N__36823));
    InMux I__8978 (
            .O(N__36860),
            .I(N__36823));
    InMux I__8977 (
            .O(N__36859),
            .I(N__36823));
    InMux I__8976 (
            .O(N__36858),
            .I(N__36823));
    InMux I__8975 (
            .O(N__36855),
            .I(N__36818));
    InMux I__8974 (
            .O(N__36854),
            .I(N__36818));
    LocalMux I__8973 (
            .O(N__36851),
            .I(N__36813));
    LocalMux I__8972 (
            .O(N__36848),
            .I(N__36813));
    Span4Mux_v I__8971 (
            .O(N__36845),
            .I(N__36809));
    InMux I__8970 (
            .O(N__36844),
            .I(N__36803));
    InMux I__8969 (
            .O(N__36841),
            .I(N__36803));
    LocalMux I__8968 (
            .O(N__36838),
            .I(N__36800));
    LocalMux I__8967 (
            .O(N__36835),
            .I(N__36797));
    LocalMux I__8966 (
            .O(N__36832),
            .I(N__36790));
    LocalMux I__8965 (
            .O(N__36823),
            .I(N__36790));
    LocalMux I__8964 (
            .O(N__36818),
            .I(N__36790));
    Span4Mux_s3_h I__8963 (
            .O(N__36813),
            .I(N__36787));
    InMux I__8962 (
            .O(N__36812),
            .I(N__36784));
    Span4Mux_h I__8961 (
            .O(N__36809),
            .I(N__36781));
    InMux I__8960 (
            .O(N__36808),
            .I(N__36778));
    LocalMux I__8959 (
            .O(N__36803),
            .I(N__36773));
    Sp12to4 I__8958 (
            .O(N__36800),
            .I(N__36773));
    Span4Mux_s3_v I__8957 (
            .O(N__36797),
            .I(N__36770));
    Span4Mux_s3_v I__8956 (
            .O(N__36790),
            .I(N__36767));
    Span4Mux_h I__8955 (
            .O(N__36787),
            .I(N__36762));
    LocalMux I__8954 (
            .O(N__36784),
            .I(N__36762));
    Span4Mux_h I__8953 (
            .O(N__36781),
            .I(N__36759));
    LocalMux I__8952 (
            .O(N__36778),
            .I(N__36756));
    Span12Mux_s8_h I__8951 (
            .O(N__36773),
            .I(N__36753));
    Span4Mux_h I__8950 (
            .O(N__36770),
            .I(N__36746));
    Span4Mux_h I__8949 (
            .O(N__36767),
            .I(N__36746));
    Span4Mux_v I__8948 (
            .O(N__36762),
            .I(N__36746));
    Odrv4 I__8947 (
            .O(N__36759),
            .I(\Inst_core.resetCmd ));
    Odrv12 I__8946 (
            .O(N__36756),
            .I(\Inst_core.resetCmd ));
    Odrv12 I__8945 (
            .O(N__36753),
            .I(\Inst_core.resetCmd ));
    Odrv4 I__8944 (
            .O(N__36746),
            .I(\Inst_core.resetCmd ));
    IoInMux I__8943 (
            .O(N__36737),
            .I(N__36734));
    LocalMux I__8942 (
            .O(N__36734),
            .I(debugleds_c_0));
    InMux I__8941 (
            .O(N__36731),
            .I(N__36725));
    InMux I__8940 (
            .O(N__36730),
            .I(N__36725));
    LocalMux I__8939 (
            .O(N__36725),
            .I(N__36722));
    Span12Mux_s0_h I__8938 (
            .O(N__36722),
            .I(N__36719));
    Odrv12 I__8937 (
            .O(N__36719),
            .I(busy));
    CascadeMux I__8936 (
            .O(N__36716),
            .I(N__36713));
    InMux I__8935 (
            .O(N__36713),
            .I(N__36710));
    LocalMux I__8934 (
            .O(N__36710),
            .I(\Inst_core.Inst_controller.nstate_1_N_825_0 ));
    CascadeMux I__8933 (
            .O(N__36707),
            .I(N__36702));
    InMux I__8932 (
            .O(N__36706),
            .I(N__36692));
    InMux I__8931 (
            .O(N__36705),
            .I(N__36692));
    InMux I__8930 (
            .O(N__36702),
            .I(N__36692));
    InMux I__8929 (
            .O(N__36701),
            .I(N__36692));
    LocalMux I__8928 (
            .O(N__36692),
            .I(\Inst_core.Inst_controller.n320 ));
    InMux I__8927 (
            .O(N__36689),
            .I(N__36680));
    InMux I__8926 (
            .O(N__36688),
            .I(N__36680));
    InMux I__8925 (
            .O(N__36687),
            .I(N__36680));
    LocalMux I__8924 (
            .O(N__36680),
            .I(N__36677));
    Odrv12 I__8923 (
            .O(N__36677),
            .I(\Inst_core.Inst_controller.nstate_1_N_829_0 ));
    InMux I__8922 (
            .O(N__36674),
            .I(N__36671));
    LocalMux I__8921 (
            .O(N__36671),
            .I(\Inst_core.Inst_controller.n2717 ));
    CEMux I__8920 (
            .O(N__36668),
            .I(N__36665));
    LocalMux I__8919 (
            .O(N__36665),
            .I(N__36659));
    InMux I__8918 (
            .O(N__36664),
            .I(N__36651));
    InMux I__8917 (
            .O(N__36663),
            .I(N__36651));
    CascadeMux I__8916 (
            .O(N__36662),
            .I(N__36648));
    Span4Mux_h I__8915 (
            .O(N__36659),
            .I(N__36640));
    InMux I__8914 (
            .O(N__36658),
            .I(N__36637));
    CascadeMux I__8913 (
            .O(N__36657),
            .I(N__36630));
    CascadeMux I__8912 (
            .O(N__36656),
            .I(N__36627));
    LocalMux I__8911 (
            .O(N__36651),
            .I(N__36622));
    InMux I__8910 (
            .O(N__36648),
            .I(N__36613));
    InMux I__8909 (
            .O(N__36647),
            .I(N__36613));
    InMux I__8908 (
            .O(N__36646),
            .I(N__36613));
    InMux I__8907 (
            .O(N__36645),
            .I(N__36613));
    InMux I__8906 (
            .O(N__36644),
            .I(N__36606));
    CEMux I__8905 (
            .O(N__36643),
            .I(N__36603));
    Span4Mux_v I__8904 (
            .O(N__36640),
            .I(N__36598));
    LocalMux I__8903 (
            .O(N__36637),
            .I(N__36598));
    InMux I__8902 (
            .O(N__36636),
            .I(N__36589));
    InMux I__8901 (
            .O(N__36635),
            .I(N__36589));
    InMux I__8900 (
            .O(N__36634),
            .I(N__36589));
    InMux I__8899 (
            .O(N__36633),
            .I(N__36589));
    InMux I__8898 (
            .O(N__36630),
            .I(N__36580));
    InMux I__8897 (
            .O(N__36627),
            .I(N__36580));
    InMux I__8896 (
            .O(N__36626),
            .I(N__36580));
    InMux I__8895 (
            .O(N__36625),
            .I(N__36580));
    Span4Mux_s2_v I__8894 (
            .O(N__36622),
            .I(N__36577));
    LocalMux I__8893 (
            .O(N__36613),
            .I(N__36574));
    InMux I__8892 (
            .O(N__36612),
            .I(N__36571));
    InMux I__8891 (
            .O(N__36611),
            .I(N__36566));
    InMux I__8890 (
            .O(N__36610),
            .I(N__36566));
    CEMux I__8889 (
            .O(N__36609),
            .I(N__36558));
    LocalMux I__8888 (
            .O(N__36606),
            .I(N__36554));
    LocalMux I__8887 (
            .O(N__36603),
            .I(N__36548));
    Span4Mux_h I__8886 (
            .O(N__36598),
            .I(N__36548));
    LocalMux I__8885 (
            .O(N__36589),
            .I(N__36543));
    LocalMux I__8884 (
            .O(N__36580),
            .I(N__36543));
    Span4Mux_h I__8883 (
            .O(N__36577),
            .I(N__36534));
    Span4Mux_s2_v I__8882 (
            .O(N__36574),
            .I(N__36534));
    LocalMux I__8881 (
            .O(N__36571),
            .I(N__36534));
    LocalMux I__8880 (
            .O(N__36566),
            .I(N__36534));
    InMux I__8879 (
            .O(N__36565),
            .I(N__36525));
    InMux I__8878 (
            .O(N__36564),
            .I(N__36525));
    InMux I__8877 (
            .O(N__36563),
            .I(N__36525));
    InMux I__8876 (
            .O(N__36562),
            .I(N__36525));
    CEMux I__8875 (
            .O(N__36561),
            .I(N__36522));
    LocalMux I__8874 (
            .O(N__36558),
            .I(N__36519));
    InMux I__8873 (
            .O(N__36557),
            .I(N__36516));
    Span4Mux_v I__8872 (
            .O(N__36554),
            .I(N__36513));
    CascadeMux I__8871 (
            .O(N__36553),
            .I(N__36509));
    Span4Mux_h I__8870 (
            .O(N__36548),
            .I(N__36503));
    Span4Mux_h I__8869 (
            .O(N__36543),
            .I(N__36503));
    Sp12to4 I__8868 (
            .O(N__36534),
            .I(N__36498));
    LocalMux I__8867 (
            .O(N__36525),
            .I(N__36498));
    LocalMux I__8866 (
            .O(N__36522),
            .I(N__36495));
    Span4Mux_h I__8865 (
            .O(N__36519),
            .I(N__36492));
    LocalMux I__8864 (
            .O(N__36516),
            .I(N__36489));
    Span4Mux_h I__8863 (
            .O(N__36513),
            .I(N__36486));
    InMux I__8862 (
            .O(N__36512),
            .I(N__36479));
    InMux I__8861 (
            .O(N__36509),
            .I(N__36479));
    InMux I__8860 (
            .O(N__36508),
            .I(N__36479));
    Sp12to4 I__8859 (
            .O(N__36503),
            .I(N__36474));
    Span12Mux_s1_h I__8858 (
            .O(N__36498),
            .I(N__36474));
    Span4Mux_s1_v I__8857 (
            .O(N__36495),
            .I(N__36469));
    Span4Mux_v I__8856 (
            .O(N__36492),
            .I(N__36469));
    Span4Mux_s1_h I__8855 (
            .O(N__36489),
            .I(N__36462));
    Span4Mux_h I__8854 (
            .O(N__36486),
            .I(N__36462));
    LocalMux I__8853 (
            .O(N__36479),
            .I(N__36462));
    Span12Mux_v I__8852 (
            .O(N__36474),
            .I(N__36459));
    Odrv4 I__8851 (
            .O(N__36469),
            .I(sampleReady));
    Odrv4 I__8850 (
            .O(N__36462),
            .I(sampleReady));
    Odrv12 I__8849 (
            .O(N__36459),
            .I(sampleReady));
    InMux I__8848 (
            .O(N__36452),
            .I(N__36438));
    InMux I__8847 (
            .O(N__36451),
            .I(N__36438));
    InMux I__8846 (
            .O(N__36450),
            .I(N__36438));
    InMux I__8845 (
            .O(N__36449),
            .I(N__36438));
    InMux I__8844 (
            .O(N__36448),
            .I(N__36433));
    InMux I__8843 (
            .O(N__36447),
            .I(N__36433));
    LocalMux I__8842 (
            .O(N__36438),
            .I(\Inst_core.n318 ));
    LocalMux I__8841 (
            .O(N__36433),
            .I(\Inst_core.n318 ));
    CascadeMux I__8840 (
            .O(N__36428),
            .I(\Inst_core.Inst_controller.n2717_cascade_ ));
    InMux I__8839 (
            .O(N__36425),
            .I(N__36415));
    InMux I__8838 (
            .O(N__36424),
            .I(N__36415));
    InMux I__8837 (
            .O(N__36423),
            .I(N__36415));
    CascadeMux I__8836 (
            .O(N__36422),
            .I(N__36403));
    LocalMux I__8835 (
            .O(N__36415),
            .I(N__36396));
    InMux I__8834 (
            .O(N__36414),
            .I(N__36393));
    InMux I__8833 (
            .O(N__36413),
            .I(N__36390));
    InMux I__8832 (
            .O(N__36412),
            .I(N__36375));
    InMux I__8831 (
            .O(N__36411),
            .I(N__36375));
    InMux I__8830 (
            .O(N__36410),
            .I(N__36375));
    InMux I__8829 (
            .O(N__36409),
            .I(N__36375));
    InMux I__8828 (
            .O(N__36408),
            .I(N__36375));
    InMux I__8827 (
            .O(N__36407),
            .I(N__36375));
    InMux I__8826 (
            .O(N__36406),
            .I(N__36375));
    InMux I__8825 (
            .O(N__36403),
            .I(N__36370));
    InMux I__8824 (
            .O(N__36402),
            .I(N__36370));
    InMux I__8823 (
            .O(N__36401),
            .I(N__36363));
    InMux I__8822 (
            .O(N__36400),
            .I(N__36363));
    InMux I__8821 (
            .O(N__36399),
            .I(N__36363));
    Span4Mux_h I__8820 (
            .O(N__36396),
            .I(N__36358));
    LocalMux I__8819 (
            .O(N__36393),
            .I(N__36358));
    LocalMux I__8818 (
            .O(N__36390),
            .I(N__36353));
    LocalMux I__8817 (
            .O(N__36375),
            .I(N__36353));
    LocalMux I__8816 (
            .O(N__36370),
            .I(N__36350));
    LocalMux I__8815 (
            .O(N__36363),
            .I(N__36347));
    Span4Mux_v I__8814 (
            .O(N__36358),
            .I(N__36343));
    Span4Mux_s2_v I__8813 (
            .O(N__36353),
            .I(N__36340));
    Span4Mux_v I__8812 (
            .O(N__36350),
            .I(N__36334));
    Span4Mux_v I__8811 (
            .O(N__36347),
            .I(N__36334));
    InMux I__8810 (
            .O(N__36346),
            .I(N__36331));
    Span4Mux_v I__8809 (
            .O(N__36343),
            .I(N__36326));
    Span4Mux_v I__8808 (
            .O(N__36340),
            .I(N__36326));
    CascadeMux I__8807 (
            .O(N__36339),
            .I(N__36322));
    Sp12to4 I__8806 (
            .O(N__36334),
            .I(N__36310));
    LocalMux I__8805 (
            .O(N__36331),
            .I(N__36310));
    Sp12to4 I__8804 (
            .O(N__36326),
            .I(N__36310));
    InMux I__8803 (
            .O(N__36325),
            .I(N__36305));
    InMux I__8802 (
            .O(N__36322),
            .I(N__36305));
    InMux I__8801 (
            .O(N__36321),
            .I(N__36298));
    InMux I__8800 (
            .O(N__36320),
            .I(N__36298));
    InMux I__8799 (
            .O(N__36319),
            .I(N__36298));
    InMux I__8798 (
            .O(N__36318),
            .I(N__36293));
    InMux I__8797 (
            .O(N__36317),
            .I(N__36293));
    Span12Mux_s11_h I__8796 (
            .O(N__36310),
            .I(N__36290));
    LocalMux I__8795 (
            .O(N__36305),
            .I(send));
    LocalMux I__8794 (
            .O(N__36298),
            .I(send));
    LocalMux I__8793 (
            .O(N__36293),
            .I(send));
    Odrv12 I__8792 (
            .O(N__36290),
            .I(send));
    InMux I__8791 (
            .O(N__36281),
            .I(N__36278));
    LocalMux I__8790 (
            .O(N__36278),
            .I(\Inst_core.Inst_controller.n2 ));
    InMux I__8789 (
            .O(N__36275),
            .I(N__36270));
    InMux I__8788 (
            .O(N__36274),
            .I(N__36265));
    InMux I__8787 (
            .O(N__36273),
            .I(N__36265));
    LocalMux I__8786 (
            .O(N__36270),
            .I(\Inst_core.Inst_controller.counter_0 ));
    LocalMux I__8785 (
            .O(N__36265),
            .I(\Inst_core.Inst_controller.counter_0 ));
    InMux I__8784 (
            .O(N__36260),
            .I(bfn_12_12_0_));
    InMux I__8783 (
            .O(N__36257),
            .I(N__36252));
    InMux I__8782 (
            .O(N__36256),
            .I(N__36249));
    InMux I__8781 (
            .O(N__36255),
            .I(N__36246));
    LocalMux I__8780 (
            .O(N__36252),
            .I(\Inst_core.Inst_controller.counter_1 ));
    LocalMux I__8779 (
            .O(N__36249),
            .I(\Inst_core.Inst_controller.counter_1 ));
    LocalMux I__8778 (
            .O(N__36246),
            .I(\Inst_core.Inst_controller.counter_1 ));
    InMux I__8777 (
            .O(N__36239),
            .I(\Inst_core.Inst_controller.n7845 ));
    InMux I__8776 (
            .O(N__36236),
            .I(N__36231));
    InMux I__8775 (
            .O(N__36235),
            .I(N__36228));
    InMux I__8774 (
            .O(N__36234),
            .I(N__36225));
    LocalMux I__8773 (
            .O(N__36231),
            .I(\Inst_core.Inst_controller.counter_2 ));
    LocalMux I__8772 (
            .O(N__36228),
            .I(\Inst_core.Inst_controller.counter_2 ));
    LocalMux I__8771 (
            .O(N__36225),
            .I(\Inst_core.Inst_controller.counter_2 ));
    InMux I__8770 (
            .O(N__36218),
            .I(\Inst_core.Inst_controller.n7846 ));
    CascadeMux I__8769 (
            .O(N__36215),
            .I(N__36212));
    InMux I__8768 (
            .O(N__36212),
            .I(N__36208));
    InMux I__8767 (
            .O(N__36211),
            .I(N__36205));
    LocalMux I__8766 (
            .O(N__36208),
            .I(N__36199));
    LocalMux I__8765 (
            .O(N__36205),
            .I(N__36199));
    InMux I__8764 (
            .O(N__36204),
            .I(N__36196));
    Span4Mux_h I__8763 (
            .O(N__36199),
            .I(N__36193));
    LocalMux I__8762 (
            .O(N__36196),
            .I(\Inst_core.Inst_controller.counter_3 ));
    Odrv4 I__8761 (
            .O(N__36193),
            .I(\Inst_core.Inst_controller.counter_3 ));
    InMux I__8760 (
            .O(N__36188),
            .I(\Inst_core.Inst_controller.n7847 ));
    InMux I__8759 (
            .O(N__36185),
            .I(N__36181));
    CascadeMux I__8758 (
            .O(N__36184),
            .I(N__36178));
    LocalMux I__8757 (
            .O(N__36181),
            .I(N__36172));
    InMux I__8756 (
            .O(N__36178),
            .I(N__36169));
    InMux I__8755 (
            .O(N__36177),
            .I(N__36162));
    InMux I__8754 (
            .O(N__36176),
            .I(N__36162));
    InMux I__8753 (
            .O(N__36175),
            .I(N__36162));
    Span4Mux_v I__8752 (
            .O(N__36172),
            .I(N__36155));
    LocalMux I__8751 (
            .O(N__36169),
            .I(N__36155));
    LocalMux I__8750 (
            .O(N__36162),
            .I(N__36152));
    InMux I__8749 (
            .O(N__36161),
            .I(N__36147));
    InMux I__8748 (
            .O(N__36160),
            .I(N__36147));
    Span4Mux_v I__8747 (
            .O(N__36155),
            .I(N__36143));
    Span4Mux_v I__8746 (
            .O(N__36152),
            .I(N__36140));
    LocalMux I__8745 (
            .O(N__36147),
            .I(N__36137));
    InMux I__8744 (
            .O(N__36146),
            .I(N__36134));
    Odrv4 I__8743 (
            .O(N__36143),
            .I(cmd_24));
    Odrv4 I__8742 (
            .O(N__36140),
            .I(cmd_24));
    Odrv4 I__8741 (
            .O(N__36137),
            .I(cmd_24));
    LocalMux I__8740 (
            .O(N__36134),
            .I(cmd_24));
    CascadeMux I__8739 (
            .O(N__36125),
            .I(N__36122));
    InMux I__8738 (
            .O(N__36122),
            .I(N__36119));
    LocalMux I__8737 (
            .O(N__36119),
            .I(N__36115));
    InMux I__8736 (
            .O(N__36118),
            .I(N__36112));
    Span4Mux_h I__8735 (
            .O(N__36115),
            .I(N__36109));
    LocalMux I__8734 (
            .O(N__36112),
            .I(configRegister_16_adj_1344));
    Odrv4 I__8733 (
            .O(N__36109),
            .I(configRegister_16_adj_1344));
    InMux I__8732 (
            .O(N__36104),
            .I(N__36100));
    InMux I__8731 (
            .O(N__36103),
            .I(N__36096));
    LocalMux I__8730 (
            .O(N__36100),
            .I(N__36093));
    InMux I__8729 (
            .O(N__36099),
            .I(N__36085));
    LocalMux I__8728 (
            .O(N__36096),
            .I(N__36080));
    Span4Mux_v I__8727 (
            .O(N__36093),
            .I(N__36080));
    InMux I__8726 (
            .O(N__36092),
            .I(N__36077));
    InMux I__8725 (
            .O(N__36091),
            .I(N__36074));
    InMux I__8724 (
            .O(N__36090),
            .I(N__36071));
    InMux I__8723 (
            .O(N__36089),
            .I(N__36068));
    InMux I__8722 (
            .O(N__36088),
            .I(N__36065));
    LocalMux I__8721 (
            .O(N__36085),
            .I(N__36062));
    Span4Mux_v I__8720 (
            .O(N__36080),
            .I(N__36057));
    LocalMux I__8719 (
            .O(N__36077),
            .I(N__36057));
    LocalMux I__8718 (
            .O(N__36074),
            .I(N__36052));
    LocalMux I__8717 (
            .O(N__36071),
            .I(N__36052));
    LocalMux I__8716 (
            .O(N__36068),
            .I(N__36047));
    LocalMux I__8715 (
            .O(N__36065),
            .I(N__36047));
    Span4Mux_h I__8714 (
            .O(N__36062),
            .I(N__36044));
    Span4Mux_s3_h I__8713 (
            .O(N__36057),
            .I(N__36041));
    Span4Mux_s3_h I__8712 (
            .O(N__36052),
            .I(N__36038));
    Span4Mux_h I__8711 (
            .O(N__36047),
            .I(N__36033));
    Span4Mux_h I__8710 (
            .O(N__36044),
            .I(N__36033));
    Span4Mux_h I__8709 (
            .O(N__36041),
            .I(N__36030));
    Span4Mux_h I__8708 (
            .O(N__36038),
            .I(N__36027));
    Odrv4 I__8707 (
            .O(N__36033),
            .I(wrtrigval_3));
    Odrv4 I__8706 (
            .O(N__36030),
            .I(wrtrigval_3));
    Odrv4 I__8705 (
            .O(N__36027),
            .I(wrtrigval_3));
    InMux I__8704 (
            .O(N__36020),
            .I(N__36017));
    LocalMux I__8703 (
            .O(N__36017),
            .I(N__36014));
    Span4Mux_s2_v I__8702 (
            .O(N__36014),
            .I(N__36011));
    Span4Mux_v I__8701 (
            .O(N__36011),
            .I(N__36007));
    InMux I__8700 (
            .O(N__36010),
            .I(N__36004));
    Odrv4 I__8699 (
            .O(N__36007),
            .I(valueRegister_0_adj_1376));
    LocalMux I__8698 (
            .O(N__36004),
            .I(valueRegister_0_adj_1376));
    InMux I__8697 (
            .O(N__35999),
            .I(N__35990));
    InMux I__8696 (
            .O(N__35998),
            .I(N__35990));
    InMux I__8695 (
            .O(N__35997),
            .I(N__35985));
    InMux I__8694 (
            .O(N__35996),
            .I(N__35981));
    InMux I__8693 (
            .O(N__35995),
            .I(N__35978));
    LocalMux I__8692 (
            .O(N__35990),
            .I(N__35975));
    InMux I__8691 (
            .O(N__35989),
            .I(N__35972));
    InMux I__8690 (
            .O(N__35988),
            .I(N__35969));
    LocalMux I__8689 (
            .O(N__35985),
            .I(N__35966));
    InMux I__8688 (
            .O(N__35984),
            .I(N__35963));
    LocalMux I__8687 (
            .O(N__35981),
            .I(N__35958));
    LocalMux I__8686 (
            .O(N__35978),
            .I(N__35958));
    Span4Mux_s2_v I__8685 (
            .O(N__35975),
            .I(N__35951));
    LocalMux I__8684 (
            .O(N__35972),
            .I(N__35948));
    LocalMux I__8683 (
            .O(N__35969),
            .I(N__35945));
    Span4Mux_v I__8682 (
            .O(N__35966),
            .I(N__35940));
    LocalMux I__8681 (
            .O(N__35963),
            .I(N__35940));
    Span4Mux_v I__8680 (
            .O(N__35958),
            .I(N__35937));
    InMux I__8679 (
            .O(N__35957),
            .I(N__35934));
    InMux I__8678 (
            .O(N__35956),
            .I(N__35929));
    InMux I__8677 (
            .O(N__35955),
            .I(N__35929));
    CascadeMux I__8676 (
            .O(N__35954),
            .I(N__35922));
    Span4Mux_v I__8675 (
            .O(N__35951),
            .I(N__35917));
    Span4Mux_v I__8674 (
            .O(N__35948),
            .I(N__35917));
    Span4Mux_v I__8673 (
            .O(N__35945),
            .I(N__35914));
    Span4Mux_v I__8672 (
            .O(N__35940),
            .I(N__35911));
    Sp12to4 I__8671 (
            .O(N__35937),
            .I(N__35904));
    LocalMux I__8670 (
            .O(N__35934),
            .I(N__35904));
    LocalMux I__8669 (
            .O(N__35929),
            .I(N__35904));
    InMux I__8668 (
            .O(N__35928),
            .I(N__35901));
    InMux I__8667 (
            .O(N__35927),
            .I(N__35896));
    InMux I__8666 (
            .O(N__35926),
            .I(N__35896));
    InMux I__8665 (
            .O(N__35925),
            .I(N__35893));
    InMux I__8664 (
            .O(N__35922),
            .I(N__35890));
    Odrv4 I__8663 (
            .O(N__35917),
            .I(cmd_8));
    Odrv4 I__8662 (
            .O(N__35914),
            .I(cmd_8));
    Odrv4 I__8661 (
            .O(N__35911),
            .I(cmd_8));
    Odrv12 I__8660 (
            .O(N__35904),
            .I(cmd_8));
    LocalMux I__8659 (
            .O(N__35901),
            .I(cmd_8));
    LocalMux I__8658 (
            .O(N__35896),
            .I(cmd_8));
    LocalMux I__8657 (
            .O(N__35893),
            .I(cmd_8));
    LocalMux I__8656 (
            .O(N__35890),
            .I(cmd_8));
    CascadeMux I__8655 (
            .O(N__35873),
            .I(N__35869));
    InMux I__8654 (
            .O(N__35872),
            .I(N__35866));
    InMux I__8653 (
            .O(N__35869),
            .I(N__35863));
    LocalMux I__8652 (
            .O(N__35866),
            .I(bwd_0));
    LocalMux I__8651 (
            .O(N__35863),
            .I(bwd_0));
    InMux I__8650 (
            .O(N__35858),
            .I(N__35845));
    InMux I__8649 (
            .O(N__35857),
            .I(N__35836));
    InMux I__8648 (
            .O(N__35856),
            .I(N__35836));
    InMux I__8647 (
            .O(N__35855),
            .I(N__35836));
    InMux I__8646 (
            .O(N__35854),
            .I(N__35836));
    InMux I__8645 (
            .O(N__35853),
            .I(N__35826));
    InMux I__8644 (
            .O(N__35852),
            .I(N__35826));
    InMux I__8643 (
            .O(N__35851),
            .I(N__35821));
    InMux I__8642 (
            .O(N__35850),
            .I(N__35821));
    InMux I__8641 (
            .O(N__35849),
            .I(N__35817));
    InMux I__8640 (
            .O(N__35848),
            .I(N__35814));
    LocalMux I__8639 (
            .O(N__35845),
            .I(N__35808));
    LocalMux I__8638 (
            .O(N__35836),
            .I(N__35808));
    InMux I__8637 (
            .O(N__35835),
            .I(N__35803));
    InMux I__8636 (
            .O(N__35834),
            .I(N__35803));
    InMux I__8635 (
            .O(N__35833),
            .I(N__35796));
    InMux I__8634 (
            .O(N__35832),
            .I(N__35791));
    InMux I__8633 (
            .O(N__35831),
            .I(N__35787));
    LocalMux I__8632 (
            .O(N__35826),
            .I(N__35782));
    LocalMux I__8631 (
            .O(N__35821),
            .I(N__35782));
    InMux I__8630 (
            .O(N__35820),
            .I(N__35779));
    LocalMux I__8629 (
            .O(N__35817),
            .I(N__35774));
    LocalMux I__8628 (
            .O(N__35814),
            .I(N__35774));
    InMux I__8627 (
            .O(N__35813),
            .I(N__35771));
    Span4Mux_v I__8626 (
            .O(N__35808),
            .I(N__35766));
    LocalMux I__8625 (
            .O(N__35803),
            .I(N__35766));
    InMux I__8624 (
            .O(N__35802),
            .I(N__35763));
    InMux I__8623 (
            .O(N__35801),
            .I(N__35758));
    InMux I__8622 (
            .O(N__35800),
            .I(N__35758));
    InMux I__8621 (
            .O(N__35799),
            .I(N__35755));
    LocalMux I__8620 (
            .O(N__35796),
            .I(N__35752));
    InMux I__8619 (
            .O(N__35795),
            .I(N__35749));
    InMux I__8618 (
            .O(N__35794),
            .I(N__35746));
    LocalMux I__8617 (
            .O(N__35791),
            .I(N__35743));
    InMux I__8616 (
            .O(N__35790),
            .I(N__35740));
    LocalMux I__8615 (
            .O(N__35787),
            .I(N__35733));
    Span4Mux_v I__8614 (
            .O(N__35782),
            .I(N__35733));
    LocalMux I__8613 (
            .O(N__35779),
            .I(N__35733));
    Span4Mux_v I__8612 (
            .O(N__35774),
            .I(N__35730));
    LocalMux I__8611 (
            .O(N__35771),
            .I(N__35725));
    Span4Mux_v I__8610 (
            .O(N__35766),
            .I(N__35725));
    LocalMux I__8609 (
            .O(N__35763),
            .I(N__35720));
    LocalMux I__8608 (
            .O(N__35758),
            .I(N__35720));
    LocalMux I__8607 (
            .O(N__35755),
            .I(N__35715));
    Span4Mux_s3_v I__8606 (
            .O(N__35752),
            .I(N__35715));
    LocalMux I__8605 (
            .O(N__35749),
            .I(N__35708));
    LocalMux I__8604 (
            .O(N__35746),
            .I(N__35708));
    Span4Mux_v I__8603 (
            .O(N__35743),
            .I(N__35708));
    LocalMux I__8602 (
            .O(N__35740),
            .I(N__35701));
    Span4Mux_v I__8601 (
            .O(N__35733),
            .I(N__35701));
    Span4Mux_h I__8600 (
            .O(N__35730),
            .I(N__35701));
    Span4Mux_h I__8599 (
            .O(N__35725),
            .I(N__35698));
    Span4Mux_s3_v I__8598 (
            .O(N__35720),
            .I(N__35691));
    Span4Mux_h I__8597 (
            .O(N__35715),
            .I(N__35691));
    Span4Mux_v I__8596 (
            .O(N__35708),
            .I(N__35691));
    Span4Mux_h I__8595 (
            .O(N__35701),
            .I(N__35688));
    Odrv4 I__8594 (
            .O(N__35698),
            .I(wrtrigcfg_2));
    Odrv4 I__8593 (
            .O(N__35691),
            .I(wrtrigcfg_2));
    Odrv4 I__8592 (
            .O(N__35688),
            .I(wrtrigcfg_2));
    InMux I__8591 (
            .O(N__35681),
            .I(N__35677));
    InMux I__8590 (
            .O(N__35680),
            .I(N__35673));
    LocalMux I__8589 (
            .O(N__35677),
            .I(N__35668));
    InMux I__8588 (
            .O(N__35676),
            .I(N__35665));
    LocalMux I__8587 (
            .O(N__35673),
            .I(N__35662));
    InMux I__8586 (
            .O(N__35672),
            .I(N__35659));
    InMux I__8585 (
            .O(N__35671),
            .I(N__35656));
    Span4Mux_s1_h I__8584 (
            .O(N__35668),
            .I(N__35651));
    LocalMux I__8583 (
            .O(N__35665),
            .I(N__35651));
    Span4Mux_v I__8582 (
            .O(N__35662),
            .I(N__35644));
    LocalMux I__8581 (
            .O(N__35659),
            .I(N__35644));
    LocalMux I__8580 (
            .O(N__35656),
            .I(N__35644));
    Span4Mux_v I__8579 (
            .O(N__35651),
            .I(N__35640));
    Span4Mux_v I__8578 (
            .O(N__35644),
            .I(N__35637));
    InMux I__8577 (
            .O(N__35643),
            .I(N__35634));
    Span4Mux_h I__8576 (
            .O(N__35640),
            .I(N__35630));
    Span4Mux_h I__8575 (
            .O(N__35637),
            .I(N__35627));
    LocalMux I__8574 (
            .O(N__35634),
            .I(N__35624));
    InMux I__8573 (
            .O(N__35633),
            .I(N__35621));
    Odrv4 I__8572 (
            .O(N__35630),
            .I(cmd_34));
    Odrv4 I__8571 (
            .O(N__35627),
            .I(cmd_34));
    Odrv12 I__8570 (
            .O(N__35624),
            .I(cmd_34));
    LocalMux I__8569 (
            .O(N__35621),
            .I(cmd_34));
    InMux I__8568 (
            .O(N__35612),
            .I(N__35607));
    CascadeMux I__8567 (
            .O(N__35611),
            .I(N__35602));
    CascadeMux I__8566 (
            .O(N__35610),
            .I(N__35597));
    LocalMux I__8565 (
            .O(N__35607),
            .I(N__35594));
    InMux I__8564 (
            .O(N__35606),
            .I(N__35591));
    CascadeMux I__8563 (
            .O(N__35605),
            .I(N__35588));
    InMux I__8562 (
            .O(N__35602),
            .I(N__35585));
    InMux I__8561 (
            .O(N__35601),
            .I(N__35582));
    CascadeMux I__8560 (
            .O(N__35600),
            .I(N__35579));
    InMux I__8559 (
            .O(N__35597),
            .I(N__35575));
    Span4Mux_h I__8558 (
            .O(N__35594),
            .I(N__35570));
    LocalMux I__8557 (
            .O(N__35591),
            .I(N__35570));
    InMux I__8556 (
            .O(N__35588),
            .I(N__35567));
    LocalMux I__8555 (
            .O(N__35585),
            .I(N__35562));
    LocalMux I__8554 (
            .O(N__35582),
            .I(N__35562));
    InMux I__8553 (
            .O(N__35579),
            .I(N__35559));
    CascadeMux I__8552 (
            .O(N__35578),
            .I(N__35556));
    LocalMux I__8551 (
            .O(N__35575),
            .I(N__35553));
    Span4Mux_h I__8550 (
            .O(N__35570),
            .I(N__35548));
    LocalMux I__8549 (
            .O(N__35567),
            .I(N__35548));
    Span4Mux_s3_v I__8548 (
            .O(N__35562),
            .I(N__35543));
    LocalMux I__8547 (
            .O(N__35559),
            .I(N__35543));
    InMux I__8546 (
            .O(N__35556),
            .I(N__35540));
    Span4Mux_v I__8545 (
            .O(N__35553),
            .I(N__35536));
    Span4Mux_s3_v I__8544 (
            .O(N__35548),
            .I(N__35529));
    Span4Mux_h I__8543 (
            .O(N__35543),
            .I(N__35529));
    LocalMux I__8542 (
            .O(N__35540),
            .I(N__35529));
    InMux I__8541 (
            .O(N__35539),
            .I(N__35526));
    Odrv4 I__8540 (
            .O(N__35536),
            .I(configRegister_26_adj_1337));
    Odrv4 I__8539 (
            .O(N__35529),
            .I(configRegister_26_adj_1337));
    LocalMux I__8538 (
            .O(N__35526),
            .I(configRegister_26_adj_1337));
    InMux I__8537 (
            .O(N__35519),
            .I(N__35500));
    InMux I__8536 (
            .O(N__35518),
            .I(N__35500));
    InMux I__8535 (
            .O(N__35517),
            .I(N__35497));
    InMux I__8534 (
            .O(N__35516),
            .I(N__35492));
    InMux I__8533 (
            .O(N__35515),
            .I(N__35492));
    InMux I__8532 (
            .O(N__35514),
            .I(N__35479));
    InMux I__8531 (
            .O(N__35513),
            .I(N__35479));
    InMux I__8530 (
            .O(N__35512),
            .I(N__35479));
    InMux I__8529 (
            .O(N__35511),
            .I(N__35479));
    InMux I__8528 (
            .O(N__35510),
            .I(N__35479));
    InMux I__8527 (
            .O(N__35509),
            .I(N__35479));
    InMux I__8526 (
            .O(N__35508),
            .I(N__35473));
    InMux I__8525 (
            .O(N__35507),
            .I(N__35470));
    InMux I__8524 (
            .O(N__35506),
            .I(N__35467));
    InMux I__8523 (
            .O(N__35505),
            .I(N__35462));
    LocalMux I__8522 (
            .O(N__35500),
            .I(N__35453));
    LocalMux I__8521 (
            .O(N__35497),
            .I(N__35453));
    LocalMux I__8520 (
            .O(N__35492),
            .I(N__35453));
    LocalMux I__8519 (
            .O(N__35479),
            .I(N__35453));
    InMux I__8518 (
            .O(N__35478),
            .I(N__35448));
    InMux I__8517 (
            .O(N__35477),
            .I(N__35448));
    InMux I__8516 (
            .O(N__35476),
            .I(N__35445));
    LocalMux I__8515 (
            .O(N__35473),
            .I(N__35434));
    LocalMux I__8514 (
            .O(N__35470),
            .I(N__35434));
    LocalMux I__8513 (
            .O(N__35467),
            .I(N__35434));
    InMux I__8512 (
            .O(N__35466),
            .I(N__35427));
    InMux I__8511 (
            .O(N__35465),
            .I(N__35427));
    LocalMux I__8510 (
            .O(N__35462),
            .I(N__35422));
    Span4Mux_v I__8509 (
            .O(N__35453),
            .I(N__35422));
    LocalMux I__8508 (
            .O(N__35448),
            .I(N__35417));
    LocalMux I__8507 (
            .O(N__35445),
            .I(N__35417));
    InMux I__8506 (
            .O(N__35444),
            .I(N__35414));
    InMux I__8505 (
            .O(N__35443),
            .I(N__35411));
    InMux I__8504 (
            .O(N__35442),
            .I(N__35408));
    CascadeMux I__8503 (
            .O(N__35441),
            .I(N__35402));
    Span4Mux_v I__8502 (
            .O(N__35434),
            .I(N__35398));
    InMux I__8501 (
            .O(N__35433),
            .I(N__35395));
    InMux I__8500 (
            .O(N__35432),
            .I(N__35392));
    LocalMux I__8499 (
            .O(N__35427),
            .I(N__35383));
    Span4Mux_s3_h I__8498 (
            .O(N__35422),
            .I(N__35383));
    Span4Mux_h I__8497 (
            .O(N__35417),
            .I(N__35383));
    LocalMux I__8496 (
            .O(N__35414),
            .I(N__35383));
    LocalMux I__8495 (
            .O(N__35411),
            .I(N__35378));
    LocalMux I__8494 (
            .O(N__35408),
            .I(N__35378));
    InMux I__8493 (
            .O(N__35407),
            .I(N__35375));
    InMux I__8492 (
            .O(N__35406),
            .I(N__35366));
    InMux I__8491 (
            .O(N__35405),
            .I(N__35366));
    InMux I__8490 (
            .O(N__35402),
            .I(N__35366));
    InMux I__8489 (
            .O(N__35401),
            .I(N__35366));
    Span4Mux_h I__8488 (
            .O(N__35398),
            .I(N__35357));
    LocalMux I__8487 (
            .O(N__35395),
            .I(N__35357));
    LocalMux I__8486 (
            .O(N__35392),
            .I(N__35357));
    Span4Mux_v I__8485 (
            .O(N__35383),
            .I(N__35354));
    Span4Mux_s2_h I__8484 (
            .O(N__35378),
            .I(N__35347));
    LocalMux I__8483 (
            .O(N__35375),
            .I(N__35347));
    LocalMux I__8482 (
            .O(N__35366),
            .I(N__35347));
    InMux I__8481 (
            .O(N__35365),
            .I(N__35344));
    InMux I__8480 (
            .O(N__35364),
            .I(N__35341));
    Span4Mux_v I__8479 (
            .O(N__35357),
            .I(N__35338));
    Span4Mux_h I__8478 (
            .O(N__35354),
            .I(N__35335));
    Span4Mux_h I__8477 (
            .O(N__35347),
            .I(N__35328));
    LocalMux I__8476 (
            .O(N__35344),
            .I(N__35328));
    LocalMux I__8475 (
            .O(N__35341),
            .I(N__35328));
    Span4Mux_h I__8474 (
            .O(N__35338),
            .I(N__35325));
    Span4Mux_h I__8473 (
            .O(N__35335),
            .I(N__35322));
    Span4Mux_v I__8472 (
            .O(N__35328),
            .I(N__35319));
    Odrv4 I__8471 (
            .O(N__35325),
            .I(wrsize));
    Odrv4 I__8470 (
            .O(N__35322),
            .I(wrsize));
    Odrv4 I__8469 (
            .O(N__35319),
            .I(wrsize));
    InMux I__8468 (
            .O(N__35312),
            .I(N__35302));
    InMux I__8467 (
            .O(N__35311),
            .I(N__35302));
    InMux I__8466 (
            .O(N__35310),
            .I(N__35299));
    InMux I__8465 (
            .O(N__35309),
            .I(N__35296));
    InMux I__8464 (
            .O(N__35308),
            .I(N__35293));
    InMux I__8463 (
            .O(N__35307),
            .I(N__35290));
    LocalMux I__8462 (
            .O(N__35302),
            .I(N__35286));
    LocalMux I__8461 (
            .O(N__35299),
            .I(N__35283));
    LocalMux I__8460 (
            .O(N__35296),
            .I(N__35280));
    LocalMux I__8459 (
            .O(N__35293),
            .I(N__35277));
    LocalMux I__8458 (
            .O(N__35290),
            .I(N__35274));
    InMux I__8457 (
            .O(N__35289),
            .I(N__35271));
    Span4Mux_v I__8456 (
            .O(N__35286),
            .I(N__35267));
    Span4Mux_s2_h I__8455 (
            .O(N__35283),
            .I(N__35264));
    Span4Mux_s2_h I__8454 (
            .O(N__35280),
            .I(N__35261));
    Span4Mux_v I__8453 (
            .O(N__35277),
            .I(N__35254));
    Span4Mux_h I__8452 (
            .O(N__35274),
            .I(N__35254));
    LocalMux I__8451 (
            .O(N__35271),
            .I(N__35254));
    InMux I__8450 (
            .O(N__35270),
            .I(N__35251));
    Odrv4 I__8449 (
            .O(N__35267),
            .I(cmd_20));
    Odrv4 I__8448 (
            .O(N__35264),
            .I(cmd_20));
    Odrv4 I__8447 (
            .O(N__35261),
            .I(cmd_20));
    Odrv4 I__8446 (
            .O(N__35254),
            .I(cmd_20));
    LocalMux I__8445 (
            .O(N__35251),
            .I(cmd_20));
    CascadeMux I__8444 (
            .O(N__35240),
            .I(N__35237));
    InMux I__8443 (
            .O(N__35237),
            .I(N__35234));
    LocalMux I__8442 (
            .O(N__35234),
            .I(N__35230));
    InMux I__8441 (
            .O(N__35233),
            .I(N__35227));
    Span4Mux_v I__8440 (
            .O(N__35230),
            .I(N__35224));
    LocalMux I__8439 (
            .O(N__35227),
            .I(bwd_12));
    Odrv4 I__8438 (
            .O(N__35224),
            .I(bwd_12));
    InMux I__8437 (
            .O(N__35219),
            .I(N__35216));
    LocalMux I__8436 (
            .O(N__35216),
            .I(N__35212));
    InMux I__8435 (
            .O(N__35215),
            .I(N__35209));
    Sp12to4 I__8434 (
            .O(N__35212),
            .I(N__35204));
    LocalMux I__8433 (
            .O(N__35209),
            .I(N__35204));
    Span12Mux_v I__8432 (
            .O(N__35204),
            .I(N__35201));
    Odrv12 I__8431 (
            .O(N__35201),
            .I(\Inst_core.nstate_1_N_831_0 ));
    CascadeMux I__8430 (
            .O(N__35198),
            .I(N__35194));
    InMux I__8429 (
            .O(N__35197),
            .I(N__35189));
    InMux I__8428 (
            .O(N__35194),
            .I(N__35189));
    LocalMux I__8427 (
            .O(N__35189),
            .I(\Inst_core.Inst_controller.n321 ));
    InMux I__8426 (
            .O(N__35186),
            .I(N__35179));
    InMux I__8425 (
            .O(N__35185),
            .I(N__35179));
    InMux I__8424 (
            .O(N__35184),
            .I(N__35176));
    LocalMux I__8423 (
            .O(N__35179),
            .I(\Inst_core.Inst_controller.nstate_1_N_827_1 ));
    LocalMux I__8422 (
            .O(N__35176),
            .I(\Inst_core.Inst_controller.nstate_1_N_827_1 ));
    CascadeMux I__8421 (
            .O(N__35171),
            .I(N__35168));
    InMux I__8420 (
            .O(N__35168),
            .I(N__35164));
    InMux I__8419 (
            .O(N__35167),
            .I(N__35161));
    LocalMux I__8418 (
            .O(N__35164),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8 ));
    LocalMux I__8417 (
            .O(N__35161),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8 ));
    InMux I__8416 (
            .O(N__35156),
            .I(N__35152));
    InMux I__8415 (
            .O(N__35155),
            .I(N__35149));
    LocalMux I__8414 (
            .O(N__35152),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13 ));
    LocalMux I__8413 (
            .O(N__35149),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13 ));
    CascadeMux I__8412 (
            .O(N__35144),
            .I(N__35140));
    CascadeMux I__8411 (
            .O(N__35143),
            .I(N__35137));
    InMux I__8410 (
            .O(N__35140),
            .I(N__35134));
    InMux I__8409 (
            .O(N__35137),
            .I(N__35131));
    LocalMux I__8408 (
            .O(N__35134),
            .I(N__35128));
    LocalMux I__8407 (
            .O(N__35131),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5 ));
    Odrv4 I__8406 (
            .O(N__35128),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5 ));
    CascadeMux I__8405 (
            .O(N__35123),
            .I(N__35119));
    InMux I__8404 (
            .O(N__35122),
            .I(N__35116));
    InMux I__8403 (
            .O(N__35119),
            .I(N__35113));
    LocalMux I__8402 (
            .O(N__35116),
            .I(N__35110));
    LocalMux I__8401 (
            .O(N__35113),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3 ));
    Odrv4 I__8400 (
            .O(N__35110),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3 ));
    InMux I__8399 (
            .O(N__35105),
            .I(N__35102));
    LocalMux I__8398 (
            .O(N__35102),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n26 ));
    InMux I__8397 (
            .O(N__35099),
            .I(N__35096));
    LocalMux I__8396 (
            .O(N__35096),
            .I(N__35092));
    InMux I__8395 (
            .O(N__35095),
            .I(N__35089));
    Odrv4 I__8394 (
            .O(N__35092),
            .I(configRegister_1));
    LocalMux I__8393 (
            .O(N__35089),
            .I(configRegister_1));
    InMux I__8392 (
            .O(N__35084),
            .I(N__35080));
    InMux I__8391 (
            .O(N__35083),
            .I(N__35077));
    LocalMux I__8390 (
            .O(N__35080),
            .I(N__35074));
    LocalMux I__8389 (
            .O(N__35077),
            .I(configRegister_16));
    Odrv4 I__8388 (
            .O(N__35074),
            .I(configRegister_16));
    InMux I__8387 (
            .O(N__35069),
            .I(N__35064));
    InMux I__8386 (
            .O(N__35068),
            .I(N__35061));
    CascadeMux I__8385 (
            .O(N__35067),
            .I(N__35042));
    LocalMux I__8384 (
            .O(N__35064),
            .I(N__35037));
    LocalMux I__8383 (
            .O(N__35061),
            .I(N__35037));
    InMux I__8382 (
            .O(N__35060),
            .I(N__35034));
    InMux I__8381 (
            .O(N__35059),
            .I(N__35031));
    InMux I__8380 (
            .O(N__35058),
            .I(N__35026));
    InMux I__8379 (
            .O(N__35057),
            .I(N__35026));
    InMux I__8378 (
            .O(N__35056),
            .I(N__35023));
    InMux I__8377 (
            .O(N__35055),
            .I(N__35018));
    InMux I__8376 (
            .O(N__35054),
            .I(N__35018));
    InMux I__8375 (
            .O(N__35053),
            .I(N__35014));
    InMux I__8374 (
            .O(N__35052),
            .I(N__35011));
    InMux I__8373 (
            .O(N__35051),
            .I(N__35006));
    InMux I__8372 (
            .O(N__35050),
            .I(N__35006));
    InMux I__8371 (
            .O(N__35049),
            .I(N__34997));
    InMux I__8370 (
            .O(N__35048),
            .I(N__34997));
    InMux I__8369 (
            .O(N__35047),
            .I(N__34997));
    InMux I__8368 (
            .O(N__35046),
            .I(N__34997));
    InMux I__8367 (
            .O(N__35045),
            .I(N__34992));
    InMux I__8366 (
            .O(N__35042),
            .I(N__34989));
    Span4Mux_v I__8365 (
            .O(N__35037),
            .I(N__34980));
    LocalMux I__8364 (
            .O(N__35034),
            .I(N__34980));
    LocalMux I__8363 (
            .O(N__35031),
            .I(N__34980));
    LocalMux I__8362 (
            .O(N__35026),
            .I(N__34980));
    LocalMux I__8361 (
            .O(N__35023),
            .I(N__34977));
    LocalMux I__8360 (
            .O(N__35018),
            .I(N__34974));
    InMux I__8359 (
            .O(N__35017),
            .I(N__34971));
    LocalMux I__8358 (
            .O(N__35014),
            .I(N__34966));
    LocalMux I__8357 (
            .O(N__35011),
            .I(N__34966));
    LocalMux I__8356 (
            .O(N__35006),
            .I(N__34955));
    LocalMux I__8355 (
            .O(N__34997),
            .I(N__34952));
    InMux I__8354 (
            .O(N__34996),
            .I(N__34947));
    InMux I__8353 (
            .O(N__34995),
            .I(N__34947));
    LocalMux I__8352 (
            .O(N__34992),
            .I(N__34944));
    LocalMux I__8351 (
            .O(N__34989),
            .I(N__34941));
    Span4Mux_h I__8350 (
            .O(N__34980),
            .I(N__34936));
    Span4Mux_h I__8349 (
            .O(N__34977),
            .I(N__34936));
    Span4Mux_h I__8348 (
            .O(N__34974),
            .I(N__34929));
    LocalMux I__8347 (
            .O(N__34971),
            .I(N__34929));
    Span4Mux_h I__8346 (
            .O(N__34966),
            .I(N__34926));
    InMux I__8345 (
            .O(N__34965),
            .I(N__34923));
    InMux I__8344 (
            .O(N__34964),
            .I(N__34920));
    InMux I__8343 (
            .O(N__34963),
            .I(N__34911));
    InMux I__8342 (
            .O(N__34962),
            .I(N__34911));
    InMux I__8341 (
            .O(N__34961),
            .I(N__34911));
    InMux I__8340 (
            .O(N__34960),
            .I(N__34911));
    InMux I__8339 (
            .O(N__34959),
            .I(N__34906));
    InMux I__8338 (
            .O(N__34958),
            .I(N__34906));
    Span4Mux_v I__8337 (
            .O(N__34955),
            .I(N__34901));
    Span4Mux_v I__8336 (
            .O(N__34952),
            .I(N__34901));
    LocalMux I__8335 (
            .O(N__34947),
            .I(N__34898));
    Span4Mux_h I__8334 (
            .O(N__34944),
            .I(N__34891));
    Span4Mux_h I__8333 (
            .O(N__34941),
            .I(N__34891));
    Span4Mux_v I__8332 (
            .O(N__34936),
            .I(N__34891));
    InMux I__8331 (
            .O(N__34935),
            .I(N__34886));
    InMux I__8330 (
            .O(N__34934),
            .I(N__34886));
    Span4Mux_h I__8329 (
            .O(N__34929),
            .I(N__34881));
    Span4Mux_h I__8328 (
            .O(N__34926),
            .I(N__34881));
    LocalMux I__8327 (
            .O(N__34923),
            .I(N__34870));
    LocalMux I__8326 (
            .O(N__34920),
            .I(N__34870));
    LocalMux I__8325 (
            .O(N__34911),
            .I(N__34870));
    LocalMux I__8324 (
            .O(N__34906),
            .I(N__34870));
    Sp12to4 I__8323 (
            .O(N__34901),
            .I(N__34870));
    Span4Mux_v I__8322 (
            .O(N__34898),
            .I(N__34867));
    Span4Mux_v I__8321 (
            .O(N__34891),
            .I(N__34864));
    LocalMux I__8320 (
            .O(N__34886),
            .I(N__34857));
    Sp12to4 I__8319 (
            .O(N__34881),
            .I(N__34857));
    Span12Mux_s8_h I__8318 (
            .O(N__34870),
            .I(N__34857));
    Odrv4 I__8317 (
            .O(N__34867),
            .I(n3753));
    Odrv4 I__8316 (
            .O(N__34864),
            .I(n3753));
    Odrv12 I__8315 (
            .O(N__34857),
            .I(n3753));
    CascadeMux I__8314 (
            .O(N__34850),
            .I(N__34847));
    InMux I__8313 (
            .O(N__34847),
            .I(N__34836));
    InMux I__8312 (
            .O(N__34846),
            .I(N__34827));
    InMux I__8311 (
            .O(N__34845),
            .I(N__34827));
    InMux I__8310 (
            .O(N__34844),
            .I(N__34827));
    InMux I__8309 (
            .O(N__34843),
            .I(N__34827));
    CascadeMux I__8308 (
            .O(N__34842),
            .I(N__34822));
    InMux I__8307 (
            .O(N__34841),
            .I(N__34814));
    CascadeMux I__8306 (
            .O(N__34840),
            .I(N__34811));
    CascadeMux I__8305 (
            .O(N__34839),
            .I(N__34806));
    LocalMux I__8304 (
            .O(N__34836),
            .I(N__34793));
    LocalMux I__8303 (
            .O(N__34827),
            .I(N__34790));
    CascadeMux I__8302 (
            .O(N__34826),
            .I(N__34786));
    InMux I__8301 (
            .O(N__34825),
            .I(N__34783));
    InMux I__8300 (
            .O(N__34822),
            .I(N__34778));
    InMux I__8299 (
            .O(N__34821),
            .I(N__34778));
    InMux I__8298 (
            .O(N__34820),
            .I(N__34768));
    InMux I__8297 (
            .O(N__34819),
            .I(N__34768));
    InMux I__8296 (
            .O(N__34818),
            .I(N__34763));
    InMux I__8295 (
            .O(N__34817),
            .I(N__34763));
    LocalMux I__8294 (
            .O(N__34814),
            .I(N__34760));
    InMux I__8293 (
            .O(N__34811),
            .I(N__34757));
    InMux I__8292 (
            .O(N__34810),
            .I(N__34754));
    InMux I__8291 (
            .O(N__34809),
            .I(N__34747));
    InMux I__8290 (
            .O(N__34806),
            .I(N__34747));
    InMux I__8289 (
            .O(N__34805),
            .I(N__34747));
    InMux I__8288 (
            .O(N__34804),
            .I(N__34744));
    InMux I__8287 (
            .O(N__34803),
            .I(N__34739));
    InMux I__8286 (
            .O(N__34802),
            .I(N__34739));
    InMux I__8285 (
            .O(N__34801),
            .I(N__34736));
    InMux I__8284 (
            .O(N__34800),
            .I(N__34733));
    InMux I__8283 (
            .O(N__34799),
            .I(N__34730));
    InMux I__8282 (
            .O(N__34798),
            .I(N__34725));
    InMux I__8281 (
            .O(N__34797),
            .I(N__34725));
    InMux I__8280 (
            .O(N__34796),
            .I(N__34722));
    Span4Mux_v I__8279 (
            .O(N__34793),
            .I(N__34717));
    Span4Mux_v I__8278 (
            .O(N__34790),
            .I(N__34717));
    InMux I__8277 (
            .O(N__34789),
            .I(N__34712));
    InMux I__8276 (
            .O(N__34786),
            .I(N__34712));
    LocalMux I__8275 (
            .O(N__34783),
            .I(N__34707));
    LocalMux I__8274 (
            .O(N__34778),
            .I(N__34707));
    CascadeMux I__8273 (
            .O(N__34777),
            .I(N__34703));
    InMux I__8272 (
            .O(N__34776),
            .I(N__34695));
    InMux I__8271 (
            .O(N__34775),
            .I(N__34692));
    InMux I__8270 (
            .O(N__34774),
            .I(N__34687));
    InMux I__8269 (
            .O(N__34773),
            .I(N__34687));
    LocalMux I__8268 (
            .O(N__34768),
            .I(N__34680));
    LocalMux I__8267 (
            .O(N__34763),
            .I(N__34680));
    Span4Mux_h I__8266 (
            .O(N__34760),
            .I(N__34680));
    LocalMux I__8265 (
            .O(N__34757),
            .I(N__34675));
    LocalMux I__8264 (
            .O(N__34754),
            .I(N__34675));
    LocalMux I__8263 (
            .O(N__34747),
            .I(N__34672));
    LocalMux I__8262 (
            .O(N__34744),
            .I(N__34653));
    LocalMux I__8261 (
            .O(N__34739),
            .I(N__34653));
    LocalMux I__8260 (
            .O(N__34736),
            .I(N__34653));
    LocalMux I__8259 (
            .O(N__34733),
            .I(N__34653));
    LocalMux I__8258 (
            .O(N__34730),
            .I(N__34653));
    LocalMux I__8257 (
            .O(N__34725),
            .I(N__34653));
    LocalMux I__8256 (
            .O(N__34722),
            .I(N__34653));
    Span4Mux_h I__8255 (
            .O(N__34717),
            .I(N__34653));
    LocalMux I__8254 (
            .O(N__34712),
            .I(N__34653));
    Span4Mux_s3_h I__8253 (
            .O(N__34707),
            .I(N__34650));
    InMux I__8252 (
            .O(N__34706),
            .I(N__34647));
    InMux I__8251 (
            .O(N__34703),
            .I(N__34642));
    InMux I__8250 (
            .O(N__34702),
            .I(N__34642));
    InMux I__8249 (
            .O(N__34701),
            .I(N__34633));
    InMux I__8248 (
            .O(N__34700),
            .I(N__34633));
    InMux I__8247 (
            .O(N__34699),
            .I(N__34633));
    InMux I__8246 (
            .O(N__34698),
            .I(N__34633));
    LocalMux I__8245 (
            .O(N__34695),
            .I(N__34630));
    LocalMux I__8244 (
            .O(N__34692),
            .I(N__34627));
    LocalMux I__8243 (
            .O(N__34687),
            .I(N__34622));
    Span4Mux_v I__8242 (
            .O(N__34680),
            .I(N__34622));
    Span4Mux_v I__8241 (
            .O(N__34675),
            .I(N__34615));
    Span4Mux_v I__8240 (
            .O(N__34672),
            .I(N__34615));
    Span4Mux_v I__8239 (
            .O(N__34653),
            .I(N__34615));
    Span4Mux_v I__8238 (
            .O(N__34650),
            .I(N__34612));
    LocalMux I__8237 (
            .O(N__34647),
            .I(n1));
    LocalMux I__8236 (
            .O(N__34642),
            .I(n1));
    LocalMux I__8235 (
            .O(N__34633),
            .I(n1));
    Odrv4 I__8234 (
            .O(N__34630),
            .I(n1));
    Odrv4 I__8233 (
            .O(N__34627),
            .I(n1));
    Odrv4 I__8232 (
            .O(N__34622),
            .I(n1));
    Odrv4 I__8231 (
            .O(N__34615),
            .I(n1));
    Odrv4 I__8230 (
            .O(N__34612),
            .I(n1));
    InMux I__8229 (
            .O(N__34595),
            .I(N__34588));
    InMux I__8228 (
            .O(N__34594),
            .I(N__34583));
    InMux I__8227 (
            .O(N__34593),
            .I(N__34583));
    InMux I__8226 (
            .O(N__34592),
            .I(N__34579));
    InMux I__8225 (
            .O(N__34591),
            .I(N__34576));
    LocalMux I__8224 (
            .O(N__34588),
            .I(N__34573));
    LocalMux I__8223 (
            .O(N__34583),
            .I(N__34570));
    InMux I__8222 (
            .O(N__34582),
            .I(N__34565));
    LocalMux I__8221 (
            .O(N__34579),
            .I(N__34562));
    LocalMux I__8220 (
            .O(N__34576),
            .I(N__34555));
    Span4Mux_h I__8219 (
            .O(N__34573),
            .I(N__34555));
    Span4Mux_s3_v I__8218 (
            .O(N__34570),
            .I(N__34555));
    InMux I__8217 (
            .O(N__34569),
            .I(N__34552));
    InMux I__8216 (
            .O(N__34568),
            .I(N__34549));
    LocalMux I__8215 (
            .O(N__34565),
            .I(N__34546));
    Span4Mux_h I__8214 (
            .O(N__34562),
            .I(N__34543));
    Span4Mux_h I__8213 (
            .O(N__34555),
            .I(N__34540));
    LocalMux I__8212 (
            .O(N__34552),
            .I(cmd_19));
    LocalMux I__8211 (
            .O(N__34549),
            .I(cmd_19));
    Odrv12 I__8210 (
            .O(N__34546),
            .I(cmd_19));
    Odrv4 I__8209 (
            .O(N__34543),
            .I(cmd_19));
    Odrv4 I__8208 (
            .O(N__34540),
            .I(cmd_19));
    InMux I__8207 (
            .O(N__34529),
            .I(N__34524));
    InMux I__8206 (
            .O(N__34528),
            .I(N__34517));
    InMux I__8205 (
            .O(N__34527),
            .I(N__34514));
    LocalMux I__8204 (
            .O(N__34524),
            .I(N__34511));
    InMux I__8203 (
            .O(N__34523),
            .I(N__34508));
    InMux I__8202 (
            .O(N__34522),
            .I(N__34505));
    InMux I__8201 (
            .O(N__34521),
            .I(N__34502));
    InMux I__8200 (
            .O(N__34520),
            .I(N__34498));
    LocalMux I__8199 (
            .O(N__34517),
            .I(N__34495));
    LocalMux I__8198 (
            .O(N__34514),
            .I(N__34486));
    Span4Mux_h I__8197 (
            .O(N__34511),
            .I(N__34486));
    LocalMux I__8196 (
            .O(N__34508),
            .I(N__34486));
    LocalMux I__8195 (
            .O(N__34505),
            .I(N__34486));
    LocalMux I__8194 (
            .O(N__34502),
            .I(N__34483));
    CascadeMux I__8193 (
            .O(N__34501),
            .I(N__34480));
    LocalMux I__8192 (
            .O(N__34498),
            .I(N__34477));
    Span4Mux_v I__8191 (
            .O(N__34495),
            .I(N__34474));
    Span4Mux_v I__8190 (
            .O(N__34486),
            .I(N__34471));
    Span4Mux_s3_h I__8189 (
            .O(N__34483),
            .I(N__34468));
    InMux I__8188 (
            .O(N__34480),
            .I(N__34465));
    Sp12to4 I__8187 (
            .O(N__34477),
            .I(N__34462));
    Span4Mux_s1_h I__8186 (
            .O(N__34474),
            .I(N__34459));
    Span4Mux_h I__8185 (
            .O(N__34471),
            .I(N__34456));
    Span4Mux_h I__8184 (
            .O(N__34468),
            .I(N__34451));
    LocalMux I__8183 (
            .O(N__34465),
            .I(N__34451));
    Span12Mux_s8_h I__8182 (
            .O(N__34462),
            .I(N__34448));
    Span4Mux_h I__8181 (
            .O(N__34459),
            .I(N__34443));
    Span4Mux_s2_h I__8180 (
            .O(N__34456),
            .I(N__34443));
    Span4Mux_v I__8179 (
            .O(N__34451),
            .I(N__34440));
    Odrv12 I__8178 (
            .O(N__34448),
            .I(wrtrigval_1));
    Odrv4 I__8177 (
            .O(N__34443),
            .I(wrtrigval_1));
    Odrv4 I__8176 (
            .O(N__34440),
            .I(wrtrigval_1));
    InMux I__8175 (
            .O(N__34433),
            .I(N__34425));
    InMux I__8174 (
            .O(N__34432),
            .I(N__34417));
    InMux I__8173 (
            .O(N__34431),
            .I(N__34414));
    InMux I__8172 (
            .O(N__34430),
            .I(N__34411));
    CascadeMux I__8171 (
            .O(N__34429),
            .I(N__34405));
    InMux I__8170 (
            .O(N__34428),
            .I(N__34401));
    LocalMux I__8169 (
            .O(N__34425),
            .I(N__34398));
    InMux I__8168 (
            .O(N__34424),
            .I(N__34395));
    InMux I__8167 (
            .O(N__34423),
            .I(N__34392));
    InMux I__8166 (
            .O(N__34422),
            .I(N__34389));
    InMux I__8165 (
            .O(N__34421),
            .I(N__34386));
    InMux I__8164 (
            .O(N__34420),
            .I(N__34383));
    LocalMux I__8163 (
            .O(N__34417),
            .I(N__34376));
    LocalMux I__8162 (
            .O(N__34414),
            .I(N__34376));
    LocalMux I__8161 (
            .O(N__34411),
            .I(N__34376));
    InMux I__8160 (
            .O(N__34410),
            .I(N__34373));
    InMux I__8159 (
            .O(N__34409),
            .I(N__34368));
    InMux I__8158 (
            .O(N__34408),
            .I(N__34368));
    InMux I__8157 (
            .O(N__34405),
            .I(N__34363));
    InMux I__8156 (
            .O(N__34404),
            .I(N__34363));
    LocalMux I__8155 (
            .O(N__34401),
            .I(N__34360));
    Span4Mux_v I__8154 (
            .O(N__34398),
            .I(N__34357));
    LocalMux I__8153 (
            .O(N__34395),
            .I(N__34353));
    LocalMux I__8152 (
            .O(N__34392),
            .I(N__34348));
    LocalMux I__8151 (
            .O(N__34389),
            .I(N__34348));
    LocalMux I__8150 (
            .O(N__34386),
            .I(N__34341));
    LocalMux I__8149 (
            .O(N__34383),
            .I(N__34341));
    Span4Mux_v I__8148 (
            .O(N__34376),
            .I(N__34341));
    LocalMux I__8147 (
            .O(N__34373),
            .I(N__34338));
    LocalMux I__8146 (
            .O(N__34368),
            .I(N__34335));
    LocalMux I__8145 (
            .O(N__34363),
            .I(N__34332));
    Span4Mux_v I__8144 (
            .O(N__34360),
            .I(N__34327));
    Span4Mux_s2_h I__8143 (
            .O(N__34357),
            .I(N__34327));
    InMux I__8142 (
            .O(N__34356),
            .I(N__34324));
    Span4Mux_v I__8141 (
            .O(N__34353),
            .I(N__34317));
    Span4Mux_v I__8140 (
            .O(N__34348),
            .I(N__34317));
    Span4Mux_h I__8139 (
            .O(N__34341),
            .I(N__34317));
    Span4Mux_h I__8138 (
            .O(N__34338),
            .I(N__34308));
    Span4Mux_v I__8137 (
            .O(N__34335),
            .I(N__34308));
    Span4Mux_v I__8136 (
            .O(N__34332),
            .I(N__34308));
    Span4Mux_h I__8135 (
            .O(N__34327),
            .I(N__34308));
    LocalMux I__8134 (
            .O(N__34324),
            .I(cmd_14));
    Odrv4 I__8133 (
            .O(N__34317),
            .I(cmd_14));
    Odrv4 I__8132 (
            .O(N__34308),
            .I(cmd_14));
    InMux I__8131 (
            .O(N__34301),
            .I(N__34298));
    LocalMux I__8130 (
            .O(N__34298),
            .I(N__34295));
    Span4Mux_v I__8129 (
            .O(N__34295),
            .I(N__34291));
    InMux I__8128 (
            .O(N__34294),
            .I(N__34288));
    Odrv4 I__8127 (
            .O(N__34291),
            .I(valueRegister_6_adj_1290));
    LocalMux I__8126 (
            .O(N__34288),
            .I(valueRegister_6_adj_1290));
    InMux I__8125 (
            .O(N__34283),
            .I(N__34280));
    LocalMux I__8124 (
            .O(N__34280),
            .I(N__34276));
    InMux I__8123 (
            .O(N__34279),
            .I(N__34273));
    Odrv4 I__8122 (
            .O(N__34276),
            .I(configRegister_12));
    LocalMux I__8121 (
            .O(N__34273),
            .I(configRegister_12));
    InMux I__8120 (
            .O(N__34268),
            .I(N__34263));
    InMux I__8119 (
            .O(N__34267),
            .I(N__34252));
    InMux I__8118 (
            .O(N__34266),
            .I(N__34252));
    LocalMux I__8117 (
            .O(N__34263),
            .I(N__34249));
    InMux I__8116 (
            .O(N__34262),
            .I(N__34246));
    InMux I__8115 (
            .O(N__34261),
            .I(N__34241));
    InMux I__8114 (
            .O(N__34260),
            .I(N__34241));
    InMux I__8113 (
            .O(N__34259),
            .I(N__34238));
    InMux I__8112 (
            .O(N__34258),
            .I(N__34232));
    InMux I__8111 (
            .O(N__34257),
            .I(N__34232));
    LocalMux I__8110 (
            .O(N__34252),
            .I(N__34228));
    Span4Mux_s2_v I__8109 (
            .O(N__34249),
            .I(N__34223));
    LocalMux I__8108 (
            .O(N__34246),
            .I(N__34216));
    LocalMux I__8107 (
            .O(N__34241),
            .I(N__34216));
    LocalMux I__8106 (
            .O(N__34238),
            .I(N__34216));
    InMux I__8105 (
            .O(N__34237),
            .I(N__34213));
    LocalMux I__8104 (
            .O(N__34232),
            .I(N__34210));
    InMux I__8103 (
            .O(N__34231),
            .I(N__34207));
    Span4Mux_s1_v I__8102 (
            .O(N__34228),
            .I(N__34202));
    InMux I__8101 (
            .O(N__34227),
            .I(N__34197));
    InMux I__8100 (
            .O(N__34226),
            .I(N__34197));
    Span4Mux_v I__8099 (
            .O(N__34223),
            .I(N__34191));
    Span4Mux_v I__8098 (
            .O(N__34216),
            .I(N__34191));
    LocalMux I__8097 (
            .O(N__34213),
            .I(N__34188));
    Span4Mux_v I__8096 (
            .O(N__34210),
            .I(N__34183));
    LocalMux I__8095 (
            .O(N__34207),
            .I(N__34183));
    InMux I__8094 (
            .O(N__34206),
            .I(N__34180));
    CascadeMux I__8093 (
            .O(N__34205),
            .I(N__34176));
    Span4Mux_v I__8092 (
            .O(N__34202),
            .I(N__34171));
    LocalMux I__8091 (
            .O(N__34197),
            .I(N__34171));
    InMux I__8090 (
            .O(N__34196),
            .I(N__34168));
    Span4Mux_h I__8089 (
            .O(N__34191),
            .I(N__34159));
    Span4Mux_v I__8088 (
            .O(N__34188),
            .I(N__34159));
    Span4Mux_v I__8087 (
            .O(N__34183),
            .I(N__34159));
    LocalMux I__8086 (
            .O(N__34180),
            .I(N__34159));
    InMux I__8085 (
            .O(N__34179),
            .I(N__34156));
    InMux I__8084 (
            .O(N__34176),
            .I(N__34153));
    Odrv4 I__8083 (
            .O(N__34171),
            .I(cmd_9));
    LocalMux I__8082 (
            .O(N__34168),
            .I(cmd_9));
    Odrv4 I__8081 (
            .O(N__34159),
            .I(cmd_9));
    LocalMux I__8080 (
            .O(N__34156),
            .I(cmd_9));
    LocalMux I__8079 (
            .O(N__34153),
            .I(cmd_9));
    InMux I__8078 (
            .O(N__34142),
            .I(N__34139));
    LocalMux I__8077 (
            .O(N__34139),
            .I(N__34135));
    InMux I__8076 (
            .O(N__34138),
            .I(N__34132));
    Span4Mux_h I__8075 (
            .O(N__34135),
            .I(N__34129));
    LocalMux I__8074 (
            .O(N__34132),
            .I(bwd_1));
    Odrv4 I__8073 (
            .O(N__34129),
            .I(bwd_1));
    CascadeMux I__8072 (
            .O(N__34124),
            .I(N__34116));
    InMux I__8071 (
            .O(N__34123),
            .I(N__34108));
    InMux I__8070 (
            .O(N__34122),
            .I(N__34108));
    InMux I__8069 (
            .O(N__34121),
            .I(N__34092));
    InMux I__8068 (
            .O(N__34120),
            .I(N__34089));
    CascadeMux I__8067 (
            .O(N__34119),
            .I(N__34086));
    InMux I__8066 (
            .O(N__34116),
            .I(N__34075));
    InMux I__8065 (
            .O(N__34115),
            .I(N__34075));
    InMux I__8064 (
            .O(N__34114),
            .I(N__34075));
    InMux I__8063 (
            .O(N__34113),
            .I(N__34075));
    LocalMux I__8062 (
            .O(N__34108),
            .I(N__34072));
    InMux I__8061 (
            .O(N__34107),
            .I(N__34067));
    InMux I__8060 (
            .O(N__34106),
            .I(N__34067));
    InMux I__8059 (
            .O(N__34105),
            .I(N__34064));
    InMux I__8058 (
            .O(N__34104),
            .I(N__34057));
    InMux I__8057 (
            .O(N__34103),
            .I(N__34057));
    InMux I__8056 (
            .O(N__34102),
            .I(N__34057));
    InMux I__8055 (
            .O(N__34101),
            .I(N__34050));
    InMux I__8054 (
            .O(N__34100),
            .I(N__34050));
    InMux I__8053 (
            .O(N__34099),
            .I(N__34050));
    CascadeMux I__8052 (
            .O(N__34098),
            .I(N__34047));
    InMux I__8051 (
            .O(N__34097),
            .I(N__34041));
    InMux I__8050 (
            .O(N__34096),
            .I(N__34041));
    InMux I__8049 (
            .O(N__34095),
            .I(N__34038));
    LocalMux I__8048 (
            .O(N__34092),
            .I(N__34035));
    LocalMux I__8047 (
            .O(N__34089),
            .I(N__34032));
    InMux I__8046 (
            .O(N__34086),
            .I(N__34029));
    InMux I__8045 (
            .O(N__34085),
            .I(N__34026));
    InMux I__8044 (
            .O(N__34084),
            .I(N__34023));
    LocalMux I__8043 (
            .O(N__34075),
            .I(N__34020));
    Span4Mux_h I__8042 (
            .O(N__34072),
            .I(N__34015));
    LocalMux I__8041 (
            .O(N__34067),
            .I(N__34015));
    LocalMux I__8040 (
            .O(N__34064),
            .I(N__34012));
    LocalMux I__8039 (
            .O(N__34057),
            .I(N__34007));
    LocalMux I__8038 (
            .O(N__34050),
            .I(N__34007));
    InMux I__8037 (
            .O(N__34047),
            .I(N__34002));
    InMux I__8036 (
            .O(N__34046),
            .I(N__34002));
    LocalMux I__8035 (
            .O(N__34041),
            .I(N__33999));
    LocalMux I__8034 (
            .O(N__34038),
            .I(N__33988));
    Span4Mux_h I__8033 (
            .O(N__34035),
            .I(N__33988));
    Span4Mux_v I__8032 (
            .O(N__34032),
            .I(N__33988));
    LocalMux I__8031 (
            .O(N__34029),
            .I(N__33988));
    LocalMux I__8030 (
            .O(N__34026),
            .I(N__33988));
    LocalMux I__8029 (
            .O(N__34023),
            .I(N__33985));
    Span4Mux_s0_h I__8028 (
            .O(N__34020),
            .I(N__33982));
    Span4Mux_v I__8027 (
            .O(N__34015),
            .I(N__33979));
    Span4Mux_v I__8026 (
            .O(N__34012),
            .I(N__33974));
    Span4Mux_v I__8025 (
            .O(N__34007),
            .I(N__33974));
    LocalMux I__8024 (
            .O(N__34002),
            .I(N__33971));
    Span4Mux_s3_h I__8023 (
            .O(N__33999),
            .I(N__33968));
    Span4Mux_v I__8022 (
            .O(N__33988),
            .I(N__33961));
    Span4Mux_v I__8021 (
            .O(N__33985),
            .I(N__33961));
    Span4Mux_h I__8020 (
            .O(N__33982),
            .I(N__33961));
    Span4Mux_v I__8019 (
            .O(N__33979),
            .I(N__33956));
    Span4Mux_h I__8018 (
            .O(N__33974),
            .I(N__33956));
    Span4Mux_v I__8017 (
            .O(N__33971),
            .I(N__33951));
    Span4Mux_h I__8016 (
            .O(N__33968),
            .I(N__33951));
    Span4Mux_h I__8015 (
            .O(N__33961),
            .I(N__33948));
    Odrv4 I__8014 (
            .O(N__33956),
            .I(wrtrigcfg_0));
    Odrv4 I__8013 (
            .O(N__33951),
            .I(wrtrigcfg_0));
    Odrv4 I__8012 (
            .O(N__33948),
            .I(wrtrigcfg_0));
    CascadeMux I__8011 (
            .O(N__33941),
            .I(N__33937));
    InMux I__8010 (
            .O(N__33940),
            .I(N__33932));
    InMux I__8009 (
            .O(N__33937),
            .I(N__33929));
    InMux I__8008 (
            .O(N__33936),
            .I(N__33923));
    InMux I__8007 (
            .O(N__33935),
            .I(N__33923));
    LocalMux I__8006 (
            .O(N__33932),
            .I(N__33918));
    LocalMux I__8005 (
            .O(N__33929),
            .I(N__33918));
    InMux I__8004 (
            .O(N__33928),
            .I(N__33915));
    LocalMux I__8003 (
            .O(N__33923),
            .I(N__33908));
    Span4Mux_v I__8002 (
            .O(N__33918),
            .I(N__33908));
    LocalMux I__8001 (
            .O(N__33915),
            .I(N__33905));
    InMux I__8000 (
            .O(N__33914),
            .I(N__33902));
    InMux I__7999 (
            .O(N__33913),
            .I(N__33899));
    Span4Mux_h I__7998 (
            .O(N__33908),
            .I(N__33893));
    Span4Mux_v I__7997 (
            .O(N__33905),
            .I(N__33893));
    LocalMux I__7996 (
            .O(N__33902),
            .I(N__33888));
    LocalMux I__7995 (
            .O(N__33899),
            .I(N__33888));
    InMux I__7994 (
            .O(N__33898),
            .I(N__33885));
    Odrv4 I__7993 (
            .O(N__33893),
            .I(cmd_23));
    Odrv12 I__7992 (
            .O(N__33888),
            .I(cmd_23));
    LocalMux I__7991 (
            .O(N__33885),
            .I(cmd_23));
    InMux I__7990 (
            .O(N__33878),
            .I(N__33875));
    LocalMux I__7989 (
            .O(N__33875),
            .I(N__33871));
    InMux I__7988 (
            .O(N__33874),
            .I(N__33868));
    Odrv4 I__7987 (
            .O(N__33871),
            .I(configRegister_15));
    LocalMux I__7986 (
            .O(N__33868),
            .I(configRegister_15));
    CascadeMux I__7985 (
            .O(N__33863),
            .I(N__33860));
    InMux I__7984 (
            .O(N__33860),
            .I(N__33856));
    InMux I__7983 (
            .O(N__33859),
            .I(N__33853));
    LocalMux I__7982 (
            .O(N__33856),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12 ));
    LocalMux I__7981 (
            .O(N__33853),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12 ));
    InMux I__7980 (
            .O(N__33848),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7880 ));
    InMux I__7979 (
            .O(N__33845),
            .I(N__33842));
    LocalMux I__7978 (
            .O(N__33842),
            .I(N__33839));
    Span4Mux_s0_h I__7977 (
            .O(N__33839),
            .I(N__33836));
    Span4Mux_h I__7976 (
            .O(N__33836),
            .I(N__33832));
    InMux I__7975 (
            .O(N__33835),
            .I(N__33829));
    Odrv4 I__7974 (
            .O(N__33832),
            .I(configRegister_13));
    LocalMux I__7973 (
            .O(N__33829),
            .I(configRegister_13));
    InMux I__7972 (
            .O(N__33824),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7881 ));
    InMux I__7971 (
            .O(N__33821),
            .I(N__33818));
    LocalMux I__7970 (
            .O(N__33818),
            .I(N__33815));
    Span4Mux_s0_h I__7969 (
            .O(N__33815),
            .I(N__33811));
    InMux I__7968 (
            .O(N__33814),
            .I(N__33808));
    Odrv4 I__7967 (
            .O(N__33811),
            .I(configRegister_14));
    LocalMux I__7966 (
            .O(N__33808),
            .I(configRegister_14));
    CascadeMux I__7965 (
            .O(N__33803),
            .I(N__33800));
    InMux I__7964 (
            .O(N__33800),
            .I(N__33796));
    InMux I__7963 (
            .O(N__33799),
            .I(N__33793));
    LocalMux I__7962 (
            .O(N__33796),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14 ));
    LocalMux I__7961 (
            .O(N__33793),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14 ));
    InMux I__7960 (
            .O(N__33788),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7882 ));
    CascadeMux I__7959 (
            .O(N__33785),
            .I(N__33775));
    CascadeMux I__7958 (
            .O(N__33784),
            .I(N__33771));
    CascadeMux I__7957 (
            .O(N__33783),
            .I(N__33767));
    CascadeMux I__7956 (
            .O(N__33782),
            .I(N__33762));
    CascadeMux I__7955 (
            .O(N__33781),
            .I(N__33758));
    CascadeMux I__7954 (
            .O(N__33780),
            .I(N__33754));
    InMux I__7953 (
            .O(N__33779),
            .I(N__33736));
    InMux I__7952 (
            .O(N__33778),
            .I(N__33736));
    InMux I__7951 (
            .O(N__33775),
            .I(N__33736));
    InMux I__7950 (
            .O(N__33774),
            .I(N__33736));
    InMux I__7949 (
            .O(N__33771),
            .I(N__33736));
    InMux I__7948 (
            .O(N__33770),
            .I(N__33736));
    InMux I__7947 (
            .O(N__33767),
            .I(N__33736));
    InMux I__7946 (
            .O(N__33766),
            .I(N__33736));
    InMux I__7945 (
            .O(N__33765),
            .I(N__33721));
    InMux I__7944 (
            .O(N__33762),
            .I(N__33721));
    InMux I__7943 (
            .O(N__33761),
            .I(N__33721));
    InMux I__7942 (
            .O(N__33758),
            .I(N__33721));
    InMux I__7941 (
            .O(N__33757),
            .I(N__33721));
    InMux I__7940 (
            .O(N__33754),
            .I(N__33721));
    InMux I__7939 (
            .O(N__33753),
            .I(N__33721));
    LocalMux I__7938 (
            .O(N__33736),
            .I(N__33716));
    LocalMux I__7937 (
            .O(N__33721),
            .I(N__33716));
    Odrv4 I__7936 (
            .O(N__33716),
            .I(\Inst_core.n1705 ));
    InMux I__7935 (
            .O(N__33713),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7883 ));
    CascadeMux I__7934 (
            .O(N__33710),
            .I(N__33706));
    CascadeMux I__7933 (
            .O(N__33709),
            .I(N__33703));
    InMux I__7932 (
            .O(N__33706),
            .I(N__33700));
    InMux I__7931 (
            .O(N__33703),
            .I(N__33697));
    LocalMux I__7930 (
            .O(N__33700),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15 ));
    LocalMux I__7929 (
            .O(N__33697),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15 ));
    CEMux I__7928 (
            .O(N__33692),
            .I(N__33688));
    CEMux I__7927 (
            .O(N__33691),
            .I(N__33685));
    LocalMux I__7926 (
            .O(N__33688),
            .I(N__33682));
    LocalMux I__7925 (
            .O(N__33685),
            .I(N__33679));
    Span4Mux_s0_h I__7924 (
            .O(N__33682),
            .I(N__33676));
    Span4Mux_s0_h I__7923 (
            .O(N__33679),
            .I(N__33673));
    Odrv4 I__7922 (
            .O(N__33676),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4044 ));
    Odrv4 I__7921 (
            .O(N__33673),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4044 ));
    InMux I__7920 (
            .O(N__33668),
            .I(N__33665));
    LocalMux I__7919 (
            .O(N__33665),
            .I(N__33661));
    InMux I__7918 (
            .O(N__33664),
            .I(N__33658));
    Odrv4 I__7917 (
            .O(N__33661),
            .I(valueRegister_1_adj_1375));
    LocalMux I__7916 (
            .O(N__33658),
            .I(valueRegister_1_adj_1375));
    InMux I__7915 (
            .O(N__33653),
            .I(N__33648));
    CascadeMux I__7914 (
            .O(N__33652),
            .I(N__33642));
    InMux I__7913 (
            .O(N__33651),
            .I(N__33639));
    LocalMux I__7912 (
            .O(N__33648),
            .I(N__33635));
    InMux I__7911 (
            .O(N__33647),
            .I(N__33630));
    InMux I__7910 (
            .O(N__33646),
            .I(N__33627));
    CascadeMux I__7909 (
            .O(N__33645),
            .I(N__33624));
    InMux I__7908 (
            .O(N__33642),
            .I(N__33621));
    LocalMux I__7907 (
            .O(N__33639),
            .I(N__33618));
    InMux I__7906 (
            .O(N__33638),
            .I(N__33615));
    Span4Mux_v I__7905 (
            .O(N__33635),
            .I(N__33612));
    InMux I__7904 (
            .O(N__33634),
            .I(N__33609));
    InMux I__7903 (
            .O(N__33633),
            .I(N__33605));
    LocalMux I__7902 (
            .O(N__33630),
            .I(N__33602));
    LocalMux I__7901 (
            .O(N__33627),
            .I(N__33599));
    InMux I__7900 (
            .O(N__33624),
            .I(N__33596));
    LocalMux I__7899 (
            .O(N__33621),
            .I(N__33585));
    Span4Mux_v I__7898 (
            .O(N__33618),
            .I(N__33585));
    LocalMux I__7897 (
            .O(N__33615),
            .I(N__33585));
    Span4Mux_s3_h I__7896 (
            .O(N__33612),
            .I(N__33585));
    LocalMux I__7895 (
            .O(N__33609),
            .I(N__33585));
    InMux I__7894 (
            .O(N__33608),
            .I(N__33582));
    LocalMux I__7893 (
            .O(N__33605),
            .I(N__33577));
    Span12Mux_s4_h I__7892 (
            .O(N__33602),
            .I(N__33577));
    Span12Mux_s11_v I__7891 (
            .O(N__33599),
            .I(N__33574));
    LocalMux I__7890 (
            .O(N__33596),
            .I(N__33569));
    Span4Mux_h I__7889 (
            .O(N__33585),
            .I(N__33569));
    LocalMux I__7888 (
            .O(N__33582),
            .I(memoryOut_1));
    Odrv12 I__7887 (
            .O(N__33577),
            .I(memoryOut_1));
    Odrv12 I__7886 (
            .O(N__33574),
            .I(memoryOut_1));
    Odrv4 I__7885 (
            .O(N__33569),
            .I(memoryOut_1));
    CascadeMux I__7884 (
            .O(N__33560),
            .I(N__33553));
    InMux I__7883 (
            .O(N__33559),
            .I(N__33548));
    InMux I__7882 (
            .O(N__33558),
            .I(N__33545));
    CascadeMux I__7881 (
            .O(N__33557),
            .I(N__33542));
    InMux I__7880 (
            .O(N__33556),
            .I(N__33539));
    InMux I__7879 (
            .O(N__33553),
            .I(N__33535));
    InMux I__7878 (
            .O(N__33552),
            .I(N__33532));
    InMux I__7877 (
            .O(N__33551),
            .I(N__33529));
    LocalMux I__7876 (
            .O(N__33548),
            .I(N__33524));
    LocalMux I__7875 (
            .O(N__33545),
            .I(N__33524));
    InMux I__7874 (
            .O(N__33542),
            .I(N__33521));
    LocalMux I__7873 (
            .O(N__33539),
            .I(N__33518));
    InMux I__7872 (
            .O(N__33538),
            .I(N__33515));
    LocalMux I__7871 (
            .O(N__33535),
            .I(N__33511));
    LocalMux I__7870 (
            .O(N__33532),
            .I(N__33508));
    LocalMux I__7869 (
            .O(N__33529),
            .I(N__33505));
    Span4Mux_v I__7868 (
            .O(N__33524),
            .I(N__33502));
    LocalMux I__7867 (
            .O(N__33521),
            .I(N__33495));
    Span4Mux_h I__7866 (
            .O(N__33518),
            .I(N__33495));
    LocalMux I__7865 (
            .O(N__33515),
            .I(N__33495));
    InMux I__7864 (
            .O(N__33514),
            .I(N__33492));
    Span4Mux_s3_h I__7863 (
            .O(N__33511),
            .I(N__33489));
    Span12Mux_s6_v I__7862 (
            .O(N__33508),
            .I(N__33486));
    Span4Mux_h I__7861 (
            .O(N__33505),
            .I(N__33481));
    Span4Mux_h I__7860 (
            .O(N__33502),
            .I(N__33481));
    Span4Mux_s2_v I__7859 (
            .O(N__33495),
            .I(N__33478));
    LocalMux I__7858 (
            .O(N__33492),
            .I(configRegister_26_adj_1377));
    Odrv4 I__7857 (
            .O(N__33489),
            .I(configRegister_26_adj_1377));
    Odrv12 I__7856 (
            .O(N__33486),
            .I(configRegister_26_adj_1377));
    Odrv4 I__7855 (
            .O(N__33481),
            .I(configRegister_26_adj_1377));
    Odrv4 I__7854 (
            .O(N__33478),
            .I(configRegister_26_adj_1377));
    InMux I__7853 (
            .O(N__33467),
            .I(N__33464));
    LocalMux I__7852 (
            .O(N__33464),
            .I(N__33461));
    Span4Mux_s0_h I__7851 (
            .O(N__33461),
            .I(N__33458));
    Span4Mux_h I__7850 (
            .O(N__33458),
            .I(N__33453));
    InMux I__7849 (
            .O(N__33457),
            .I(N__33448));
    InMux I__7848 (
            .O(N__33456),
            .I(N__33448));
    Odrv4 I__7847 (
            .O(N__33453),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1 ));
    LocalMux I__7846 (
            .O(N__33448),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1 ));
    InMux I__7845 (
            .O(N__33443),
            .I(N__33440));
    LocalMux I__7844 (
            .O(N__33440),
            .I(N__33437));
    Span4Mux_s0_h I__7843 (
            .O(N__33437),
            .I(N__33434));
    Odrv4 I__7842 (
            .O(N__33434),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_1 ));
    SRMux I__7841 (
            .O(N__33431),
            .I(N__33428));
    LocalMux I__7840 (
            .O(N__33428),
            .I(N__33425));
    Span4Mux_s1_h I__7839 (
            .O(N__33425),
            .I(N__33422));
    Odrv4 I__7838 (
            .O(N__33422),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4760 ));
    InMux I__7837 (
            .O(N__33419),
            .I(N__33416));
    LocalMux I__7836 (
            .O(N__33416),
            .I(N__33413));
    Span4Mux_v I__7835 (
            .O(N__33413),
            .I(N__33410));
    Span4Mux_h I__7834 (
            .O(N__33410),
            .I(N__33407));
    Odrv4 I__7833 (
            .O(N__33407),
            .I(\Inst_core.Inst_trigger.stageMatch_2 ));
    InMux I__7832 (
            .O(N__33404),
            .I(N__33401));
    LocalMux I__7831 (
            .O(N__33401),
            .I(N__33398));
    Span4Mux_v I__7830 (
            .O(N__33398),
            .I(N__33395));
    Odrv4 I__7829 (
            .O(N__33395),
            .I(\Inst_core.Inst_trigger.stageMatch_3 ));
    CascadeMux I__7828 (
            .O(N__33392),
            .I(N__33389));
    InMux I__7827 (
            .O(N__33389),
            .I(N__33386));
    LocalMux I__7826 (
            .O(N__33386),
            .I(N__33383));
    Span4Mux_v I__7825 (
            .O(N__33383),
            .I(N__33380));
    Odrv4 I__7824 (
            .O(N__33380),
            .I(\Inst_core.Inst_trigger.stageMatch_1 ));
    InMux I__7823 (
            .O(N__33377),
            .I(N__33374));
    LocalMux I__7822 (
            .O(N__33374),
            .I(N__33371));
    Odrv12 I__7821 (
            .O(N__33371),
            .I(\Inst_core.Inst_trigger.stageMatch_0 ));
    CascadeMux I__7820 (
            .O(N__33368),
            .I(N__33365));
    InMux I__7819 (
            .O(N__33365),
            .I(N__33359));
    InMux I__7818 (
            .O(N__33364),
            .I(N__33359));
    LocalMux I__7817 (
            .O(N__33359),
            .I(N__33356));
    Odrv12 I__7816 (
            .O(N__33356),
            .I(\Inst_core.Inst_trigger.levelReg_1__N_590 ));
    InMux I__7815 (
            .O(N__33353),
            .I(N__33349));
    InMux I__7814 (
            .O(N__33352),
            .I(N__33346));
    LocalMux I__7813 (
            .O(N__33349),
            .I(N__33343));
    LocalMux I__7812 (
            .O(N__33346),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6 ));
    Odrv12 I__7811 (
            .O(N__33343),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6 ));
    CascadeMux I__7810 (
            .O(N__33338),
            .I(N__33334));
    InMux I__7809 (
            .O(N__33337),
            .I(N__33331));
    InMux I__7808 (
            .O(N__33334),
            .I(N__33328));
    LocalMux I__7807 (
            .O(N__33331),
            .I(N__33325));
    LocalMux I__7806 (
            .O(N__33328),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1 ));
    Odrv4 I__7805 (
            .O(N__33325),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1 ));
    CascadeMux I__7804 (
            .O(N__33320),
            .I(N__33317));
    InMux I__7803 (
            .O(N__33317),
            .I(N__33313));
    InMux I__7802 (
            .O(N__33316),
            .I(N__33310));
    LocalMux I__7801 (
            .O(N__33313),
            .I(N__33307));
    LocalMux I__7800 (
            .O(N__33310),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4 ));
    Odrv12 I__7799 (
            .O(N__33307),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4 ));
    CascadeMux I__7798 (
            .O(N__33302),
            .I(N__33298));
    InMux I__7797 (
            .O(N__33301),
            .I(N__33295));
    InMux I__7796 (
            .O(N__33298),
            .I(N__33292));
    LocalMux I__7795 (
            .O(N__33295),
            .I(N__33289));
    LocalMux I__7794 (
            .O(N__33292),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0 ));
    Odrv4 I__7793 (
            .O(N__33289),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0 ));
    InMux I__7792 (
            .O(N__33284),
            .I(N__33281));
    LocalMux I__7791 (
            .O(N__33281),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n28 ));
    CascadeMux I__7790 (
            .O(N__33278),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n25_cascade_ ));
    InMux I__7789 (
            .O(N__33275),
            .I(N__33272));
    LocalMux I__7788 (
            .O(N__33272),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n27 ));
    InMux I__7787 (
            .O(N__33269),
            .I(N__33261));
    InMux I__7786 (
            .O(N__33268),
            .I(N__33261));
    InMux I__7785 (
            .O(N__33267),
            .I(N__33253));
    InMux I__7784 (
            .O(N__33266),
            .I(N__33253));
    LocalMux I__7783 (
            .O(N__33261),
            .I(N__33250));
    InMux I__7782 (
            .O(N__33260),
            .I(N__33243));
    InMux I__7781 (
            .O(N__33259),
            .I(N__33243));
    InMux I__7780 (
            .O(N__33258),
            .I(N__33243));
    LocalMux I__7779 (
            .O(N__33253),
            .I(N__33240));
    Span4Mux_h I__7778 (
            .O(N__33250),
            .I(N__33237));
    LocalMux I__7777 (
            .O(N__33243),
            .I(N__33234));
    Span4Mux_v I__7776 (
            .O(N__33240),
            .I(N__33231));
    Odrv4 I__7775 (
            .O(N__33237),
            .I(\Inst_core.n31_adj_1132 ));
    Odrv12 I__7774 (
            .O(N__33234),
            .I(\Inst_core.n31_adj_1132 ));
    Odrv4 I__7773 (
            .O(N__33231),
            .I(\Inst_core.n31_adj_1132 ));
    InMux I__7772 (
            .O(N__33224),
            .I(N__33221));
    LocalMux I__7771 (
            .O(N__33221),
            .I(N__33217));
    InMux I__7770 (
            .O(N__33220),
            .I(N__33214));
    Odrv4 I__7769 (
            .O(N__33217),
            .I(configRegister_4));
    LocalMux I__7768 (
            .O(N__33214),
            .I(configRegister_4));
    InMux I__7767 (
            .O(N__33209),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7872 ));
    InMux I__7766 (
            .O(N__33206),
            .I(N__33203));
    LocalMux I__7765 (
            .O(N__33203),
            .I(N__33199));
    InMux I__7764 (
            .O(N__33202),
            .I(N__33196));
    Odrv4 I__7763 (
            .O(N__33199),
            .I(configRegister_5));
    LocalMux I__7762 (
            .O(N__33196),
            .I(configRegister_5));
    InMux I__7761 (
            .O(N__33191),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7873 ));
    InMux I__7760 (
            .O(N__33188),
            .I(N__33185));
    LocalMux I__7759 (
            .O(N__33185),
            .I(N__33181));
    InMux I__7758 (
            .O(N__33184),
            .I(N__33178));
    Odrv4 I__7757 (
            .O(N__33181),
            .I(configRegister_6));
    LocalMux I__7756 (
            .O(N__33178),
            .I(configRegister_6));
    InMux I__7755 (
            .O(N__33173),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7874 ));
    InMux I__7754 (
            .O(N__33170),
            .I(N__33167));
    LocalMux I__7753 (
            .O(N__33167),
            .I(N__33164));
    Span4Mux_v I__7752 (
            .O(N__33164),
            .I(N__33160));
    InMux I__7751 (
            .O(N__33163),
            .I(N__33157));
    Odrv4 I__7750 (
            .O(N__33160),
            .I(configRegister_7));
    LocalMux I__7749 (
            .O(N__33157),
            .I(configRegister_7));
    CascadeMux I__7748 (
            .O(N__33152),
            .I(N__33148));
    CascadeMux I__7747 (
            .O(N__33151),
            .I(N__33145));
    InMux I__7746 (
            .O(N__33148),
            .I(N__33142));
    InMux I__7745 (
            .O(N__33145),
            .I(N__33139));
    LocalMux I__7744 (
            .O(N__33142),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7 ));
    LocalMux I__7743 (
            .O(N__33139),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7 ));
    InMux I__7742 (
            .O(N__33134),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7875 ));
    InMux I__7741 (
            .O(N__33131),
            .I(N__33127));
    InMux I__7740 (
            .O(N__33130),
            .I(N__33124));
    LocalMux I__7739 (
            .O(N__33127),
            .I(N__33121));
    LocalMux I__7738 (
            .O(N__33124),
            .I(configRegister_8));
    Odrv12 I__7737 (
            .O(N__33121),
            .I(configRegister_8));
    InMux I__7736 (
            .O(N__33116),
            .I(bfn_12_6_0_));
    InMux I__7735 (
            .O(N__33113),
            .I(N__33110));
    LocalMux I__7734 (
            .O(N__33110),
            .I(N__33106));
    InMux I__7733 (
            .O(N__33109),
            .I(N__33103));
    Odrv4 I__7732 (
            .O(N__33106),
            .I(configRegister_9));
    LocalMux I__7731 (
            .O(N__33103),
            .I(configRegister_9));
    InMux I__7730 (
            .O(N__33098),
            .I(N__33094));
    InMux I__7729 (
            .O(N__33097),
            .I(N__33091));
    LocalMux I__7728 (
            .O(N__33094),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9 ));
    LocalMux I__7727 (
            .O(N__33091),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9 ));
    InMux I__7726 (
            .O(N__33086),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7877 ));
    InMux I__7725 (
            .O(N__33083),
            .I(N__33080));
    LocalMux I__7724 (
            .O(N__33080),
            .I(N__33077));
    Span4Mux_s3_h I__7723 (
            .O(N__33077),
            .I(N__33073));
    InMux I__7722 (
            .O(N__33076),
            .I(N__33070));
    Odrv4 I__7721 (
            .O(N__33073),
            .I(configRegister_10));
    LocalMux I__7720 (
            .O(N__33070),
            .I(configRegister_10));
    CascadeMux I__7719 (
            .O(N__33065),
            .I(N__33062));
    InMux I__7718 (
            .O(N__33062),
            .I(N__33058));
    InMux I__7717 (
            .O(N__33061),
            .I(N__33055));
    LocalMux I__7716 (
            .O(N__33058),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10 ));
    LocalMux I__7715 (
            .O(N__33055),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10 ));
    InMux I__7714 (
            .O(N__33050),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7878 ));
    InMux I__7713 (
            .O(N__33047),
            .I(N__33044));
    LocalMux I__7712 (
            .O(N__33044),
            .I(N__33041));
    Span4Mux_v I__7711 (
            .O(N__33041),
            .I(N__33037));
    InMux I__7710 (
            .O(N__33040),
            .I(N__33034));
    Odrv4 I__7709 (
            .O(N__33037),
            .I(configRegister_11));
    LocalMux I__7708 (
            .O(N__33034),
            .I(configRegister_11));
    InMux I__7707 (
            .O(N__33029),
            .I(N__33025));
    InMux I__7706 (
            .O(N__33028),
            .I(N__33022));
    LocalMux I__7705 (
            .O(N__33025),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11 ));
    LocalMux I__7704 (
            .O(N__33022),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11 ));
    InMux I__7703 (
            .O(N__33017),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7879 ));
    CascadeMux I__7702 (
            .O(N__33014),
            .I(N__33011));
    InMux I__7701 (
            .O(N__33011),
            .I(N__33007));
    InMux I__7700 (
            .O(N__33010),
            .I(N__33004));
    LocalMux I__7699 (
            .O(N__33007),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0 ));
    LocalMux I__7698 (
            .O(N__33004),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0 ));
    CascadeMux I__7697 (
            .O(N__32999),
            .I(N__32996));
    InMux I__7696 (
            .O(N__32996),
            .I(N__32992));
    InMux I__7695 (
            .O(N__32995),
            .I(N__32989));
    LocalMux I__7694 (
            .O(N__32992),
            .I(N__32986));
    LocalMux I__7693 (
            .O(N__32989),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4 ));
    Odrv4 I__7692 (
            .O(N__32986),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4 ));
    CascadeMux I__7691 (
            .O(N__32981),
            .I(N__32978));
    InMux I__7690 (
            .O(N__32978),
            .I(N__32974));
    InMux I__7689 (
            .O(N__32977),
            .I(N__32971));
    LocalMux I__7688 (
            .O(N__32974),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1 ));
    LocalMux I__7687 (
            .O(N__32971),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1 ));
    InMux I__7686 (
            .O(N__32966),
            .I(N__32963));
    LocalMux I__7685 (
            .O(N__32963),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n28 ));
    CascadeMux I__7684 (
            .O(N__32960),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n25_cascade_ ));
    InMux I__7683 (
            .O(N__32957),
            .I(N__32954));
    LocalMux I__7682 (
            .O(N__32954),
            .I(N__32951));
    Span4Mux_s3_v I__7681 (
            .O(N__32951),
            .I(N__32944));
    InMux I__7680 (
            .O(N__32950),
            .I(N__32935));
    InMux I__7679 (
            .O(N__32949),
            .I(N__32935));
    InMux I__7678 (
            .O(N__32948),
            .I(N__32935));
    InMux I__7677 (
            .O(N__32947),
            .I(N__32935));
    Odrv4 I__7676 (
            .O(N__32944),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n31 ));
    LocalMux I__7675 (
            .O(N__32935),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n31 ));
    CascadeMux I__7674 (
            .O(N__32930),
            .I(N__32926));
    InMux I__7673 (
            .O(N__32929),
            .I(N__32923));
    InMux I__7672 (
            .O(N__32926),
            .I(N__32920));
    LocalMux I__7671 (
            .O(N__32923),
            .I(N__32917));
    LocalMux I__7670 (
            .O(N__32920),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12 ));
    Odrv4 I__7669 (
            .O(N__32917),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12 ));
    InMux I__7668 (
            .O(N__32912),
            .I(N__32909));
    LocalMux I__7667 (
            .O(N__32909),
            .I(N__32905));
    InMux I__7666 (
            .O(N__32908),
            .I(N__32902));
    Odrv4 I__7665 (
            .O(N__32905),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2 ));
    LocalMux I__7664 (
            .O(N__32902),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2 ));
    CascadeMux I__7663 (
            .O(N__32897),
            .I(N__32893));
    CascadeMux I__7662 (
            .O(N__32896),
            .I(N__32890));
    InMux I__7661 (
            .O(N__32893),
            .I(N__32887));
    InMux I__7660 (
            .O(N__32890),
            .I(N__32884));
    LocalMux I__7659 (
            .O(N__32887),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7 ));
    LocalMux I__7658 (
            .O(N__32884),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7 ));
    CascadeMux I__7657 (
            .O(N__32879),
            .I(N__32876));
    InMux I__7656 (
            .O(N__32876),
            .I(N__32872));
    InMux I__7655 (
            .O(N__32875),
            .I(N__32869));
    LocalMux I__7654 (
            .O(N__32872),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10 ));
    LocalMux I__7653 (
            .O(N__32869),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10 ));
    InMux I__7652 (
            .O(N__32864),
            .I(N__32861));
    LocalMux I__7651 (
            .O(N__32861),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n27 ));
    CascadeMux I__7650 (
            .O(N__32858),
            .I(N__32855));
    InMux I__7649 (
            .O(N__32855),
            .I(N__32851));
    InMux I__7648 (
            .O(N__32854),
            .I(N__32848));
    LocalMux I__7647 (
            .O(N__32851),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3 ));
    LocalMux I__7646 (
            .O(N__32848),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3 ));
    InMux I__7645 (
            .O(N__32843),
            .I(N__32839));
    InMux I__7644 (
            .O(N__32842),
            .I(N__32836));
    LocalMux I__7643 (
            .O(N__32839),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13 ));
    LocalMux I__7642 (
            .O(N__32836),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13 ));
    CascadeMux I__7641 (
            .O(N__32831),
            .I(N__32827));
    CascadeMux I__7640 (
            .O(N__32830),
            .I(N__32824));
    InMux I__7639 (
            .O(N__32827),
            .I(N__32821));
    InMux I__7638 (
            .O(N__32824),
            .I(N__32818));
    LocalMux I__7637 (
            .O(N__32821),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5 ));
    LocalMux I__7636 (
            .O(N__32818),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5 ));
    CascadeMux I__7635 (
            .O(N__32813),
            .I(N__32810));
    InMux I__7634 (
            .O(N__32810),
            .I(N__32806));
    InMux I__7633 (
            .O(N__32809),
            .I(N__32803));
    LocalMux I__7632 (
            .O(N__32806),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8 ));
    LocalMux I__7631 (
            .O(N__32803),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8 ));
    InMux I__7630 (
            .O(N__32798),
            .I(N__32795));
    LocalMux I__7629 (
            .O(N__32795),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n26 ));
    InMux I__7628 (
            .O(N__32792),
            .I(N__32789));
    LocalMux I__7627 (
            .O(N__32789),
            .I(N__32785));
    InMux I__7626 (
            .O(N__32788),
            .I(N__32782));
    Odrv4 I__7625 (
            .O(N__32785),
            .I(configRegister_0));
    LocalMux I__7624 (
            .O(N__32782),
            .I(configRegister_0));
    InMux I__7623 (
            .O(N__32777),
            .I(N__32774));
    LocalMux I__7622 (
            .O(N__32774),
            .I(N__32771));
    Span12Mux_s11_v I__7621 (
            .O(N__32771),
            .I(N__32768));
    Odrv12 I__7620 (
            .O(N__32768),
            .I(\Inst_core.n9053 ));
    InMux I__7619 (
            .O(N__32765),
            .I(bfn_12_5_0_));
    InMux I__7618 (
            .O(N__32762),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7869 ));
    InMux I__7617 (
            .O(N__32759),
            .I(N__32756));
    LocalMux I__7616 (
            .O(N__32756),
            .I(N__32753));
    Span4Mux_v I__7615 (
            .O(N__32753),
            .I(N__32750));
    Span4Mux_h I__7614 (
            .O(N__32750),
            .I(N__32746));
    InMux I__7613 (
            .O(N__32749),
            .I(N__32743));
    Odrv4 I__7612 (
            .O(N__32746),
            .I(configRegister_2));
    LocalMux I__7611 (
            .O(N__32743),
            .I(configRegister_2));
    InMux I__7610 (
            .O(N__32738),
            .I(N__32734));
    InMux I__7609 (
            .O(N__32737),
            .I(N__32731));
    LocalMux I__7608 (
            .O(N__32734),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2 ));
    LocalMux I__7607 (
            .O(N__32731),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2 ));
    InMux I__7606 (
            .O(N__32726),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7870 ));
    InMux I__7605 (
            .O(N__32723),
            .I(N__32720));
    LocalMux I__7604 (
            .O(N__32720),
            .I(N__32716));
    InMux I__7603 (
            .O(N__32719),
            .I(N__32713));
    Odrv12 I__7602 (
            .O(N__32716),
            .I(configRegister_3));
    LocalMux I__7601 (
            .O(N__32713),
            .I(configRegister_3));
    InMux I__7600 (
            .O(N__32708),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7871 ));
    SRMux I__7599 (
            .O(N__32705),
            .I(N__32702));
    LocalMux I__7598 (
            .O(N__32702),
            .I(N__32699));
    Span4Mux_s2_h I__7597 (
            .O(N__32699),
            .I(N__32696));
    Odrv4 I__7596 (
            .O(N__32696),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4645 ));
    InMux I__7595 (
            .O(N__32693),
            .I(N__32690));
    LocalMux I__7594 (
            .O(N__32690),
            .I(N__32687));
    Span4Mux_s1_h I__7593 (
            .O(N__32687),
            .I(N__32684));
    Odrv4 I__7592 (
            .O(N__32684),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_2 ));
    InMux I__7591 (
            .O(N__32681),
            .I(N__32678));
    LocalMux I__7590 (
            .O(N__32678),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_0 ));
    InMux I__7589 (
            .O(N__32675),
            .I(N__32672));
    LocalMux I__7588 (
            .O(N__32672),
            .I(N__32669));
    Span4Mux_h I__7587 (
            .O(N__32669),
            .I(N__32666));
    Odrv4 I__7586 (
            .O(N__32666),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7_adj_1000 ));
    InMux I__7585 (
            .O(N__32663),
            .I(N__32658));
    InMux I__7584 (
            .O(N__32662),
            .I(N__32655));
    InMux I__7583 (
            .O(N__32661),
            .I(N__32652));
    LocalMux I__7582 (
            .O(N__32658),
            .I(N__32649));
    LocalMux I__7581 (
            .O(N__32655),
            .I(\Inst_core.Inst_trigger.configRegister_27 ));
    LocalMux I__7580 (
            .O(N__32652),
            .I(\Inst_core.Inst_trigger.configRegister_27 ));
    Odrv4 I__7579 (
            .O(N__32649),
            .I(\Inst_core.Inst_trigger.configRegister_27 ));
    CascadeMux I__7578 (
            .O(N__32642),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n8521_cascade_ ));
    CEMux I__7577 (
            .O(N__32639),
            .I(N__32636));
    LocalMux I__7576 (
            .O(N__32636),
            .I(N__32633));
    Span4Mux_s3_v I__7575 (
            .O(N__32633),
            .I(N__32628));
    CEMux I__7574 (
            .O(N__32632),
            .I(N__32625));
    InMux I__7573 (
            .O(N__32631),
            .I(N__32622));
    Span4Mux_s0_h I__7572 (
            .O(N__32628),
            .I(N__32613));
    LocalMux I__7571 (
            .O(N__32625),
            .I(N__32613));
    LocalMux I__7570 (
            .O(N__32622),
            .I(N__32613));
    InMux I__7569 (
            .O(N__32621),
            .I(N__32610));
    CEMux I__7568 (
            .O(N__32620),
            .I(N__32606));
    IoSpan4Mux I__7567 (
            .O(N__32613),
            .I(N__32603));
    LocalMux I__7566 (
            .O(N__32610),
            .I(N__32599));
    CEMux I__7565 (
            .O(N__32609),
            .I(N__32596));
    LocalMux I__7564 (
            .O(N__32606),
            .I(N__32591));
    IoSpan4Mux I__7563 (
            .O(N__32603),
            .I(N__32591));
    InMux I__7562 (
            .O(N__32602),
            .I(N__32588));
    Span4Mux_s3_h I__7561 (
            .O(N__32599),
            .I(N__32585));
    LocalMux I__7560 (
            .O(N__32596),
            .I(N__32578));
    Span4Mux_s3_h I__7559 (
            .O(N__32591),
            .I(N__32578));
    LocalMux I__7558 (
            .O(N__32588),
            .I(N__32578));
    Span4Mux_v I__7557 (
            .O(N__32585),
            .I(N__32575));
    Span4Mux_h I__7556 (
            .O(N__32578),
            .I(N__32572));
    Span4Mux_v I__7555 (
            .O(N__32575),
            .I(N__32569));
    Span4Mux_v I__7554 (
            .O(N__32572),
            .I(N__32566));
    Span4Mux_h I__7553 (
            .O(N__32569),
            .I(N__32563));
    Span4Mux_v I__7552 (
            .O(N__32566),
            .I(N__32560));
    Odrv4 I__7551 (
            .O(N__32563),
            .I(\Inst_core.n3670 ));
    Odrv4 I__7550 (
            .O(N__32560),
            .I(\Inst_core.n3670 ));
    InMux I__7549 (
            .O(N__32555),
            .I(N__32552));
    LocalMux I__7548 (
            .O(N__32552),
            .I(N__32549));
    Span4Mux_s2_v I__7547 (
            .O(N__32549),
            .I(N__32546));
    Odrv4 I__7546 (
            .O(N__32546),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7 ));
    InMux I__7545 (
            .O(N__32543),
            .I(N__32537));
    InMux I__7544 (
            .O(N__32542),
            .I(N__32537));
    LocalMux I__7543 (
            .O(N__32537),
            .I(N__32534));
    Span12Mux_s3_h I__7542 (
            .O(N__32534),
            .I(N__32531));
    Odrv12 I__7541 (
            .O(N__32531),
            .I(\Inst_core.Inst_trigger.stageRun_0 ));
    InMux I__7540 (
            .O(N__32528),
            .I(N__32525));
    LocalMux I__7539 (
            .O(N__32525),
            .I(N__32521));
    InMux I__7538 (
            .O(N__32524),
            .I(N__32518));
    Span4Mux_s2_h I__7537 (
            .O(N__32521),
            .I(N__32515));
    LocalMux I__7536 (
            .O(N__32518),
            .I(\Inst_core.Inst_trigger.stageRun_3 ));
    Odrv4 I__7535 (
            .O(N__32515),
            .I(\Inst_core.Inst_trigger.stageRun_3 ));
    CascadeMux I__7534 (
            .O(N__32510),
            .I(N__32507));
    InMux I__7533 (
            .O(N__32507),
            .I(N__32504));
    LocalMux I__7532 (
            .O(N__32504),
            .I(N__32500));
    InMux I__7531 (
            .O(N__32503),
            .I(N__32497));
    Span4Mux_v I__7530 (
            .O(N__32500),
            .I(N__32494));
    LocalMux I__7529 (
            .O(N__32497),
            .I(\Inst_core.stageRun_2 ));
    Odrv4 I__7528 (
            .O(N__32494),
            .I(\Inst_core.stageRun_2 ));
    InMux I__7527 (
            .O(N__32489),
            .I(N__32485));
    InMux I__7526 (
            .O(N__32488),
            .I(N__32482));
    LocalMux I__7525 (
            .O(N__32485),
            .I(\Inst_core.stageRun_1 ));
    LocalMux I__7524 (
            .O(N__32482),
            .I(\Inst_core.stageRun_1 ));
    CascadeMux I__7523 (
            .O(N__32477),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n8753_cascade_ ));
    InMux I__7522 (
            .O(N__32474),
            .I(N__32470));
    InMux I__7521 (
            .O(N__32473),
            .I(N__32467));
    LocalMux I__7520 (
            .O(N__32470),
            .I(N__32464));
    LocalMux I__7519 (
            .O(N__32467),
            .I(N__32461));
    Span4Mux_v I__7518 (
            .O(N__32464),
            .I(N__32458));
    Span4Mux_v I__7517 (
            .O(N__32461),
            .I(N__32455));
    Odrv4 I__7516 (
            .O(N__32458),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n461 ));
    Odrv4 I__7515 (
            .O(N__32455),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n461 ));
    InMux I__7514 (
            .O(N__32450),
            .I(N__32444));
    InMux I__7513 (
            .O(N__32449),
            .I(N__32444));
    LocalMux I__7512 (
            .O(N__32444),
            .I(N__32441));
    Span4Mux_s2_h I__7511 (
            .O(N__32441),
            .I(N__32435));
    InMux I__7510 (
            .O(N__32440),
            .I(N__32430));
    InMux I__7509 (
            .O(N__32439),
            .I(N__32427));
    InMux I__7508 (
            .O(N__32438),
            .I(N__32424));
    Span4Mux_v I__7507 (
            .O(N__32435),
            .I(N__32421));
    InMux I__7506 (
            .O(N__32434),
            .I(N__32416));
    InMux I__7505 (
            .O(N__32433),
            .I(N__32416));
    LocalMux I__7504 (
            .O(N__32430),
            .I(N__32413));
    LocalMux I__7503 (
            .O(N__32427),
            .I(N__32408));
    LocalMux I__7502 (
            .O(N__32424),
            .I(N__32408));
    Span4Mux_v I__7501 (
            .O(N__32421),
            .I(N__32405));
    LocalMux I__7500 (
            .O(N__32416),
            .I(\Inst_core.state_1 ));
    Odrv12 I__7499 (
            .O(N__32413),
            .I(\Inst_core.state_1 ));
    Odrv12 I__7498 (
            .O(N__32408),
            .I(\Inst_core.state_1 ));
    Odrv4 I__7497 (
            .O(N__32405),
            .I(\Inst_core.state_1 ));
    InMux I__7496 (
            .O(N__32396),
            .I(N__32393));
    LocalMux I__7495 (
            .O(N__32393),
            .I(N__32389));
    InMux I__7494 (
            .O(N__32392),
            .I(N__32386));
    Odrv12 I__7493 (
            .O(N__32389),
            .I(valueRegister_3_adj_1373));
    LocalMux I__7492 (
            .O(N__32386),
            .I(valueRegister_3_adj_1373));
    InMux I__7491 (
            .O(N__32381),
            .I(N__32378));
    LocalMux I__7490 (
            .O(N__32378),
            .I(N__32375));
    Span12Mux_s4_v I__7489 (
            .O(N__32375),
            .I(N__32370));
    InMux I__7488 (
            .O(N__32374),
            .I(N__32365));
    InMux I__7487 (
            .O(N__32373),
            .I(N__32365));
    Odrv12 I__7486 (
            .O(N__32370),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3 ));
    LocalMux I__7485 (
            .O(N__32365),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3 ));
    CascadeMux I__7484 (
            .O(N__32360),
            .I(N__32357));
    InMux I__7483 (
            .O(N__32357),
            .I(N__32354));
    LocalMux I__7482 (
            .O(N__32354),
            .I(N__32348));
    InMux I__7481 (
            .O(N__32353),
            .I(N__32345));
    InMux I__7480 (
            .O(N__32352),
            .I(N__32340));
    InMux I__7479 (
            .O(N__32351),
            .I(N__32334));
    Span4Mux_s3_h I__7478 (
            .O(N__32348),
            .I(N__32331));
    LocalMux I__7477 (
            .O(N__32345),
            .I(N__32328));
    InMux I__7476 (
            .O(N__32344),
            .I(N__32323));
    InMux I__7475 (
            .O(N__32343),
            .I(N__32323));
    LocalMux I__7474 (
            .O(N__32340),
            .I(N__32320));
    InMux I__7473 (
            .O(N__32339),
            .I(N__32317));
    InMux I__7472 (
            .O(N__32338),
            .I(N__32314));
    InMux I__7471 (
            .O(N__32337),
            .I(N__32310));
    LocalMux I__7470 (
            .O(N__32334),
            .I(N__32305));
    Span4Mux_v I__7469 (
            .O(N__32331),
            .I(N__32305));
    Sp12to4 I__7468 (
            .O(N__32328),
            .I(N__32300));
    LocalMux I__7467 (
            .O(N__32323),
            .I(N__32300));
    Span4Mux_s3_v I__7466 (
            .O(N__32320),
            .I(N__32297));
    LocalMux I__7465 (
            .O(N__32317),
            .I(N__32292));
    LocalMux I__7464 (
            .O(N__32314),
            .I(N__32292));
    InMux I__7463 (
            .O(N__32313),
            .I(N__32289));
    LocalMux I__7462 (
            .O(N__32310),
            .I(N__32286));
    Span4Mux_v I__7461 (
            .O(N__32305),
            .I(N__32283));
    Span12Mux_s11_v I__7460 (
            .O(N__32300),
            .I(N__32280));
    Span4Mux_h I__7459 (
            .O(N__32297),
            .I(N__32275));
    Span4Mux_h I__7458 (
            .O(N__32292),
            .I(N__32275));
    LocalMux I__7457 (
            .O(N__32289),
            .I(memoryOut_3));
    Odrv12 I__7456 (
            .O(N__32286),
            .I(memoryOut_3));
    Odrv4 I__7455 (
            .O(N__32283),
            .I(memoryOut_3));
    Odrv12 I__7454 (
            .O(N__32280),
            .I(memoryOut_3));
    Odrv4 I__7453 (
            .O(N__32275),
            .I(memoryOut_3));
    CascadeMux I__7452 (
            .O(N__32264),
            .I(N__32261));
    InMux I__7451 (
            .O(N__32261),
            .I(N__32258));
    LocalMux I__7450 (
            .O(N__32258),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_3 ));
    SRMux I__7449 (
            .O(N__32255),
            .I(N__32252));
    LocalMux I__7448 (
            .O(N__32252),
            .I(N__32249));
    Span4Mux_v I__7447 (
            .O(N__32249),
            .I(N__32246));
    Span4Mux_h I__7446 (
            .O(N__32246),
            .I(N__32243));
    Odrv4 I__7445 (
            .O(N__32243),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4762 ));
    InMux I__7444 (
            .O(N__32240),
            .I(N__32236));
    InMux I__7443 (
            .O(N__32239),
            .I(N__32233));
    LocalMux I__7442 (
            .O(N__32236),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6 ));
    LocalMux I__7441 (
            .O(N__32233),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6 ));
    CEMux I__7440 (
            .O(N__32228),
            .I(N__32225));
    LocalMux I__7439 (
            .O(N__32225),
            .I(N__32222));
    IoSpan4Mux I__7438 (
            .O(N__32222),
            .I(N__32219));
    Span4Mux_s0_h I__7437 (
            .O(N__32219),
            .I(N__32216));
    Odrv4 I__7436 (
            .O(N__32216),
            .I(\Inst_core.Inst_sampler.n8687 ));
    InMux I__7435 (
            .O(N__32213),
            .I(N__32210));
    LocalMux I__7434 (
            .O(N__32210),
            .I(N__32206));
    InMux I__7433 (
            .O(N__32209),
            .I(N__32203));
    Odrv12 I__7432 (
            .O(N__32206),
            .I(valueRegister_0_adj_1336));
    LocalMux I__7431 (
            .O(N__32203),
            .I(valueRegister_0_adj_1336));
    InMux I__7430 (
            .O(N__32198),
            .I(N__32194));
    CascadeMux I__7429 (
            .O(N__32197),
            .I(N__32191));
    LocalMux I__7428 (
            .O(N__32194),
            .I(N__32187));
    InMux I__7427 (
            .O(N__32191),
            .I(N__32182));
    InMux I__7426 (
            .O(N__32190),
            .I(N__32182));
    Odrv4 I__7425 (
            .O(N__32187),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0 ));
    LocalMux I__7424 (
            .O(N__32182),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0 ));
    SRMux I__7423 (
            .O(N__32177),
            .I(N__32174));
    LocalMux I__7422 (
            .O(N__32174),
            .I(N__32171));
    Span4Mux_v I__7421 (
            .O(N__32171),
            .I(N__32168));
    Span4Mux_s0_h I__7420 (
            .O(N__32168),
            .I(N__32165));
    Odrv4 I__7419 (
            .O(N__32165),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4643 ));
    InMux I__7418 (
            .O(N__32162),
            .I(N__32159));
    LocalMux I__7417 (
            .O(N__32159),
            .I(N__32156));
    Span4Mux_s1_v I__7416 (
            .O(N__32156),
            .I(N__32153));
    Odrv4 I__7415 (
            .O(N__32153),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_1 ));
    InMux I__7414 (
            .O(N__32150),
            .I(N__32147));
    LocalMux I__7413 (
            .O(N__32147),
            .I(N__32144));
    Odrv12 I__7412 (
            .O(N__32144),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_2 ));
    CascadeMux I__7411 (
            .O(N__32141),
            .I(N__32138));
    InMux I__7410 (
            .O(N__32138),
            .I(N__32135));
    LocalMux I__7409 (
            .O(N__32135),
            .I(N__32132));
    Odrv12 I__7408 (
            .O(N__32132),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_3 ));
    InMux I__7407 (
            .O(N__32129),
            .I(N__32126));
    LocalMux I__7406 (
            .O(N__32126),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_0 ));
    InMux I__7405 (
            .O(N__32123),
            .I(N__32120));
    LocalMux I__7404 (
            .O(N__32120),
            .I(N__32117));
    Span4Mux_h I__7403 (
            .O(N__32117),
            .I(N__32114));
    Span4Mux_v I__7402 (
            .O(N__32114),
            .I(N__32111));
    Odrv4 I__7401 (
            .O(N__32111),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7 ));
    CascadeMux I__7400 (
            .O(N__32108),
            .I(N__32105));
    InMux I__7399 (
            .O(N__32105),
            .I(N__32102));
    LocalMux I__7398 (
            .O(N__32102),
            .I(N__32098));
    InMux I__7397 (
            .O(N__32101),
            .I(N__32094));
    Span4Mux_v I__7396 (
            .O(N__32098),
            .I(N__32091));
    InMux I__7395 (
            .O(N__32097),
            .I(N__32088));
    LocalMux I__7394 (
            .O(N__32094),
            .I(divider_5));
    Odrv4 I__7393 (
            .O(N__32091),
            .I(divider_5));
    LocalMux I__7392 (
            .O(N__32088),
            .I(divider_5));
    InMux I__7391 (
            .O(N__32081),
            .I(N__32077));
    InMux I__7390 (
            .O(N__32080),
            .I(N__32073));
    LocalMux I__7389 (
            .O(N__32077),
            .I(N__32070));
    InMux I__7388 (
            .O(N__32076),
            .I(N__32067));
    LocalMux I__7387 (
            .O(N__32073),
            .I(N__32060));
    Span4Mux_v I__7386 (
            .O(N__32070),
            .I(N__32060));
    LocalMux I__7385 (
            .O(N__32067),
            .I(N__32060));
    Odrv4 I__7384 (
            .O(N__32060),
            .I(\Inst_core.Inst_sampler.counter_22 ));
    CascadeMux I__7383 (
            .O(N__32057),
            .I(N__32053));
    CascadeMux I__7382 (
            .O(N__32056),
            .I(N__32050));
    InMux I__7381 (
            .O(N__32053),
            .I(N__32047));
    InMux I__7380 (
            .O(N__32050),
            .I(N__32043));
    LocalMux I__7379 (
            .O(N__32047),
            .I(N__32040));
    InMux I__7378 (
            .O(N__32046),
            .I(N__32037));
    LocalMux I__7377 (
            .O(N__32043),
            .I(N__32032));
    Span12Mux_s5_h I__7376 (
            .O(N__32040),
            .I(N__32032));
    LocalMux I__7375 (
            .O(N__32037),
            .I(divider_22));
    Odrv12 I__7374 (
            .O(N__32032),
            .I(divider_22));
    InMux I__7373 (
            .O(N__32027),
            .I(N__32023));
    InMux I__7372 (
            .O(N__32026),
            .I(N__32020));
    LocalMux I__7371 (
            .O(N__32023),
            .I(N__32016));
    LocalMux I__7370 (
            .O(N__32020),
            .I(N__32013));
    InMux I__7369 (
            .O(N__32019),
            .I(N__32010));
    Span4Mux_s2_h I__7368 (
            .O(N__32016),
            .I(N__32007));
    Span4Mux_s2_h I__7367 (
            .O(N__32013),
            .I(N__32004));
    LocalMux I__7366 (
            .O(N__32010),
            .I(\Inst_core.Inst_sampler.counter_5 ));
    Odrv4 I__7365 (
            .O(N__32007),
            .I(\Inst_core.Inst_sampler.counter_5 ));
    Odrv4 I__7364 (
            .O(N__32004),
            .I(\Inst_core.Inst_sampler.counter_5 ));
    InMux I__7363 (
            .O(N__31997),
            .I(N__31994));
    LocalMux I__7362 (
            .O(N__31994),
            .I(\Inst_core.Inst_sampler.n34 ));
    InMux I__7361 (
            .O(N__31991),
            .I(N__31988));
    LocalMux I__7360 (
            .O(N__31988),
            .I(N__31985));
    Span4Mux_s3_h I__7359 (
            .O(N__31985),
            .I(N__31982));
    Odrv4 I__7358 (
            .O(N__31982),
            .I(\Inst_core.Inst_sampler.n44 ));
    InMux I__7357 (
            .O(N__31979),
            .I(N__31976));
    LocalMux I__7356 (
            .O(N__31976),
            .I(N__31973));
    Odrv4 I__7355 (
            .O(N__31973),
            .I(\Inst_core.Inst_sampler.n43 ));
    InMux I__7354 (
            .O(N__31970),
            .I(N__31967));
    LocalMux I__7353 (
            .O(N__31967),
            .I(\Inst_core.Inst_sampler.n45 ));
    InMux I__7352 (
            .O(N__31964),
            .I(N__31957));
    InMux I__7351 (
            .O(N__31963),
            .I(N__31950));
    InMux I__7350 (
            .O(N__31962),
            .I(N__31944));
    InMux I__7349 (
            .O(N__31961),
            .I(N__31944));
    InMux I__7348 (
            .O(N__31960),
            .I(N__31941));
    LocalMux I__7347 (
            .O(N__31957),
            .I(N__31938));
    IoInMux I__7346 (
            .O(N__31956),
            .I(N__31935));
    InMux I__7345 (
            .O(N__31955),
            .I(N__31932));
    InMux I__7344 (
            .O(N__31954),
            .I(N__31927));
    InMux I__7343 (
            .O(N__31953),
            .I(N__31927));
    LocalMux I__7342 (
            .O(N__31950),
            .I(N__31924));
    InMux I__7341 (
            .O(N__31949),
            .I(N__31921));
    LocalMux I__7340 (
            .O(N__31944),
            .I(N__31918));
    LocalMux I__7339 (
            .O(N__31941),
            .I(N__31915));
    Span4Mux_v I__7338 (
            .O(N__31938),
            .I(N__31912));
    LocalMux I__7337 (
            .O(N__31935),
            .I(N__31909));
    LocalMux I__7336 (
            .O(N__31932),
            .I(N__31904));
    LocalMux I__7335 (
            .O(N__31927),
            .I(N__31904));
    Span4Mux_v I__7334 (
            .O(N__31924),
            .I(N__31897));
    LocalMux I__7333 (
            .O(N__31921),
            .I(N__31897));
    Span4Mux_s2_v I__7332 (
            .O(N__31918),
            .I(N__31897));
    Span12Mux_s10_h I__7331 (
            .O(N__31915),
            .I(N__31892));
    Span4Mux_h I__7330 (
            .O(N__31912),
            .I(N__31889));
    Span4Mux_s1_h I__7329 (
            .O(N__31909),
            .I(N__31884));
    Span4Mux_h I__7328 (
            .O(N__31904),
            .I(N__31884));
    Span4Mux_h I__7327 (
            .O(N__31897),
            .I(N__31881));
    InMux I__7326 (
            .O(N__31896),
            .I(N__31876));
    InMux I__7325 (
            .O(N__31895),
            .I(N__31876));
    Span12Mux_v I__7324 (
            .O(N__31892),
            .I(N__31873));
    Odrv4 I__7323 (
            .O(N__31889),
            .I(ready50_N_581));
    Odrv4 I__7322 (
            .O(N__31884),
            .I(ready50_N_581));
    Odrv4 I__7321 (
            .O(N__31881),
            .I(ready50_N_581));
    LocalMux I__7320 (
            .O(N__31876),
            .I(ready50_N_581));
    Odrv12 I__7319 (
            .O(N__31873),
            .I(ready50_N_581));
    CascadeMux I__7318 (
            .O(N__31862),
            .I(N__31858));
    InMux I__7317 (
            .O(N__31861),
            .I(N__31854));
    InMux I__7316 (
            .O(N__31858),
            .I(N__31849));
    InMux I__7315 (
            .O(N__31857),
            .I(N__31849));
    LocalMux I__7314 (
            .O(N__31854),
            .I(\Inst_core.configRegister_27_adj_1196 ));
    LocalMux I__7313 (
            .O(N__31849),
            .I(\Inst_core.configRegister_27_adj_1196 ));
    SRMux I__7312 (
            .O(N__31844),
            .I(N__31841));
    LocalMux I__7311 (
            .O(N__31841),
            .I(N__31838));
    Span4Mux_s1_v I__7310 (
            .O(N__31838),
            .I(N__31835));
    Odrv4 I__7309 (
            .O(N__31835),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n8626 ));
    SRMux I__7308 (
            .O(N__31832),
            .I(N__31829));
    LocalMux I__7307 (
            .O(N__31829),
            .I(N__31826));
    Span4Mux_v I__7306 (
            .O(N__31826),
            .I(N__31823));
    Span4Mux_v I__7305 (
            .O(N__31823),
            .I(N__31820));
    Odrv4 I__7304 (
            .O(N__31820),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4 ));
    InMux I__7303 (
            .O(N__31817),
            .I(N__31813));
    InMux I__7302 (
            .O(N__31816),
            .I(N__31810));
    LocalMux I__7301 (
            .O(N__31813),
            .I(N__31805));
    LocalMux I__7300 (
            .O(N__31810),
            .I(N__31805));
    Span4Mux_v I__7299 (
            .O(N__31805),
            .I(N__31801));
    CascadeMux I__7298 (
            .O(N__31804),
            .I(N__31797));
    IoSpan4Mux I__7297 (
            .O(N__31801),
            .I(N__31791));
    InMux I__7296 (
            .O(N__31800),
            .I(N__31785));
    InMux I__7295 (
            .O(N__31797),
            .I(N__31782));
    InMux I__7294 (
            .O(N__31796),
            .I(N__31777));
    InMux I__7293 (
            .O(N__31795),
            .I(N__31777));
    InMux I__7292 (
            .O(N__31794),
            .I(N__31774));
    Span4Mux_s0_h I__7291 (
            .O(N__31791),
            .I(N__31771));
    InMux I__7290 (
            .O(N__31790),
            .I(N__31768));
    InMux I__7289 (
            .O(N__31789),
            .I(N__31765));
    CascadeMux I__7288 (
            .O(N__31788),
            .I(N__31762));
    LocalMux I__7287 (
            .O(N__31785),
            .I(N__31759));
    LocalMux I__7286 (
            .O(N__31782),
            .I(N__31756));
    LocalMux I__7285 (
            .O(N__31777),
            .I(N__31753));
    LocalMux I__7284 (
            .O(N__31774),
            .I(N__31750));
    Span4Mux_h I__7283 (
            .O(N__31771),
            .I(N__31743));
    LocalMux I__7282 (
            .O(N__31768),
            .I(N__31743));
    LocalMux I__7281 (
            .O(N__31765),
            .I(N__31743));
    InMux I__7280 (
            .O(N__31762),
            .I(N__31740));
    Span4Mux_v I__7279 (
            .O(N__31759),
            .I(N__31737));
    Span12Mux_s4_h I__7278 (
            .O(N__31756),
            .I(N__31734));
    Span4Mux_h I__7277 (
            .O(N__31753),
            .I(N__31729));
    Span4Mux_h I__7276 (
            .O(N__31750),
            .I(N__31729));
    Span4Mux_h I__7275 (
            .O(N__31743),
            .I(N__31726));
    LocalMux I__7274 (
            .O(N__31740),
            .I(memoryOut_0));
    Odrv4 I__7273 (
            .O(N__31737),
            .I(memoryOut_0));
    Odrv12 I__7272 (
            .O(N__31734),
            .I(memoryOut_0));
    Odrv4 I__7271 (
            .O(N__31729),
            .I(memoryOut_0));
    Odrv4 I__7270 (
            .O(N__31726),
            .I(memoryOut_0));
    InMux I__7269 (
            .O(N__31715),
            .I(N__31712));
    LocalMux I__7268 (
            .O(N__31712),
            .I(N__31709));
    Span4Mux_s0_h I__7267 (
            .O(N__31709),
            .I(N__31705));
    CascadeMux I__7266 (
            .O(N__31708),
            .I(N__31702));
    Span4Mux_h I__7265 (
            .O(N__31705),
            .I(N__31698));
    InMux I__7264 (
            .O(N__31702),
            .I(N__31693));
    InMux I__7263 (
            .O(N__31701),
            .I(N__31693));
    Odrv4 I__7262 (
            .O(N__31698),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0 ));
    LocalMux I__7261 (
            .O(N__31693),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0 ));
    CascadeMux I__7260 (
            .O(N__31688),
            .I(N__31684));
    InMux I__7259 (
            .O(N__31687),
            .I(N__31680));
    InMux I__7258 (
            .O(N__31684),
            .I(N__31677));
    InMux I__7257 (
            .O(N__31683),
            .I(N__31674));
    LocalMux I__7256 (
            .O(N__31680),
            .I(N__31671));
    LocalMux I__7255 (
            .O(N__31677),
            .I(N__31668));
    LocalMux I__7254 (
            .O(N__31674),
            .I(N__31663));
    Span4Mux_v I__7253 (
            .O(N__31671),
            .I(N__31663));
    Span4Mux_s2_h I__7252 (
            .O(N__31668),
            .I(N__31660));
    Odrv4 I__7251 (
            .O(N__31663),
            .I(divider_3));
    Odrv4 I__7250 (
            .O(N__31660),
            .I(divider_3));
    InMux I__7249 (
            .O(N__31655),
            .I(N__31651));
    InMux I__7248 (
            .O(N__31654),
            .I(N__31647));
    LocalMux I__7247 (
            .O(N__31651),
            .I(N__31644));
    InMux I__7246 (
            .O(N__31650),
            .I(N__31641));
    LocalMux I__7245 (
            .O(N__31647),
            .I(N__31634));
    Span4Mux_v I__7244 (
            .O(N__31644),
            .I(N__31634));
    LocalMux I__7243 (
            .O(N__31641),
            .I(N__31634));
    Odrv4 I__7242 (
            .O(N__31634),
            .I(\Inst_core.Inst_sampler.counter_6 ));
    InMux I__7241 (
            .O(N__31631),
            .I(N__31628));
    LocalMux I__7240 (
            .O(N__31628),
            .I(\Inst_core.Inst_sampler.n26 ));
    InMux I__7239 (
            .O(N__31625),
            .I(N__31622));
    LocalMux I__7238 (
            .O(N__31622),
            .I(N__31619));
    Span4Mux_v I__7237 (
            .O(N__31619),
            .I(N__31614));
    InMux I__7236 (
            .O(N__31618),
            .I(N__31609));
    InMux I__7235 (
            .O(N__31617),
            .I(N__31609));
    Odrv4 I__7234 (
            .O(N__31614),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3 ));
    LocalMux I__7233 (
            .O(N__31609),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3 ));
    InMux I__7232 (
            .O(N__31604),
            .I(N__31601));
    LocalMux I__7231 (
            .O(N__31601),
            .I(N__31598));
    Span4Mux_s3_h I__7230 (
            .O(N__31598),
            .I(N__31595));
    Span4Mux_v I__7229 (
            .O(N__31595),
            .I(N__31591));
    InMux I__7228 (
            .O(N__31594),
            .I(N__31588));
    Odrv4 I__7227 (
            .O(N__31591),
            .I(valueRegister_3_adj_1333));
    LocalMux I__7226 (
            .O(N__31588),
            .I(valueRegister_3_adj_1333));
    SRMux I__7225 (
            .O(N__31583),
            .I(N__31580));
    LocalMux I__7224 (
            .O(N__31580),
            .I(N__31577));
    Span4Mux_s2_h I__7223 (
            .O(N__31577),
            .I(N__31574));
    Span4Mux_s2_v I__7222 (
            .O(N__31574),
            .I(N__31571));
    Odrv4 I__7221 (
            .O(N__31571),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4755 ));
    InMux I__7220 (
            .O(N__31568),
            .I(N__31564));
    InMux I__7219 (
            .O(N__31567),
            .I(N__31561));
    LocalMux I__7218 (
            .O(N__31564),
            .I(N__31558));
    LocalMux I__7217 (
            .O(N__31561),
            .I(divider_0));
    Odrv12 I__7216 (
            .O(N__31558),
            .I(divider_0));
    InMux I__7215 (
            .O(N__31553),
            .I(N__31550));
    LocalMux I__7214 (
            .O(N__31550),
            .I(N__31545));
    InMux I__7213 (
            .O(N__31549),
            .I(N__31542));
    InMux I__7212 (
            .O(N__31548),
            .I(N__31539));
    Span4Mux_s2_h I__7211 (
            .O(N__31545),
            .I(N__31536));
    LocalMux I__7210 (
            .O(N__31542),
            .I(\Inst_core.Inst_sampler.counter_12 ));
    LocalMux I__7209 (
            .O(N__31539),
            .I(\Inst_core.Inst_sampler.counter_12 ));
    Odrv4 I__7208 (
            .O(N__31536),
            .I(\Inst_core.Inst_sampler.counter_12 ));
    CascadeMux I__7207 (
            .O(N__31529),
            .I(N__31525));
    InMux I__7206 (
            .O(N__31528),
            .I(N__31521));
    InMux I__7205 (
            .O(N__31525),
            .I(N__31518));
    InMux I__7204 (
            .O(N__31524),
            .I(N__31515));
    LocalMux I__7203 (
            .O(N__31521),
            .I(N__31510));
    LocalMux I__7202 (
            .O(N__31518),
            .I(N__31510));
    LocalMux I__7201 (
            .O(N__31515),
            .I(divider_12));
    Odrv12 I__7200 (
            .O(N__31510),
            .I(divider_12));
    InMux I__7199 (
            .O(N__31505),
            .I(N__31502));
    LocalMux I__7198 (
            .O(N__31502),
            .I(N__31499));
    Span4Mux_v I__7197 (
            .O(N__31499),
            .I(N__31494));
    InMux I__7196 (
            .O(N__31498),
            .I(N__31491));
    InMux I__7195 (
            .O(N__31497),
            .I(N__31488));
    Span4Mux_s0_h I__7194 (
            .O(N__31494),
            .I(N__31483));
    LocalMux I__7193 (
            .O(N__31491),
            .I(N__31483));
    LocalMux I__7192 (
            .O(N__31488),
            .I(\Inst_core.Inst_sampler.counter_0 ));
    Odrv4 I__7191 (
            .O(N__31483),
            .I(\Inst_core.Inst_sampler.counter_0 ));
    InMux I__7190 (
            .O(N__31478),
            .I(N__31475));
    LocalMux I__7189 (
            .O(N__31475),
            .I(\Inst_core.Inst_sampler.n25 ));
    InMux I__7188 (
            .O(N__31472),
            .I(N__31469));
    LocalMux I__7187 (
            .O(N__31469),
            .I(N__31466));
    Span4Mux_h I__7186 (
            .O(N__31466),
            .I(N__31463));
    Odrv4 I__7185 (
            .O(N__31463),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_7 ));
    InMux I__7184 (
            .O(N__31460),
            .I(N__31456));
    InMux I__7183 (
            .O(N__31459),
            .I(N__31453));
    LocalMux I__7182 (
            .O(N__31456),
            .I(N__31450));
    LocalMux I__7181 (
            .O(N__31453),
            .I(N__31447));
    Span4Mux_s3_h I__7180 (
            .O(N__31450),
            .I(N__31444));
    Span4Mux_h I__7179 (
            .O(N__31447),
            .I(N__31441));
    Odrv4 I__7178 (
            .O(N__31444),
            .I(input_c_7));
    Odrv4 I__7177 (
            .O(N__31441),
            .I(input_c_7));
    InMux I__7176 (
            .O(N__31436),
            .I(N__31432));
    CascadeMux I__7175 (
            .O(N__31435),
            .I(N__31429));
    LocalMux I__7174 (
            .O(N__31432),
            .I(N__31425));
    InMux I__7173 (
            .O(N__31429),
            .I(N__31422));
    InMux I__7172 (
            .O(N__31428),
            .I(N__31419));
    Span4Mux_h I__7171 (
            .O(N__31425),
            .I(N__31416));
    LocalMux I__7170 (
            .O(N__31422),
            .I(N__31413));
    LocalMux I__7169 (
            .O(N__31419),
            .I(\Inst_core.Inst_sync.synchronizedInput_7 ));
    Odrv4 I__7168 (
            .O(N__31416),
            .I(\Inst_core.Inst_sync.synchronizedInput_7 ));
    Odrv12 I__7167 (
            .O(N__31413),
            .I(\Inst_core.Inst_sync.synchronizedInput_7 ));
    InMux I__7166 (
            .O(N__31406),
            .I(N__31403));
    LocalMux I__7165 (
            .O(N__31403),
            .I(N__31399));
    InMux I__7164 (
            .O(N__31402),
            .I(N__31394));
    Span4Mux_v I__7163 (
            .O(N__31399),
            .I(N__31391));
    InMux I__7162 (
            .O(N__31398),
            .I(N__31388));
    CascadeMux I__7161 (
            .O(N__31397),
            .I(N__31384));
    LocalMux I__7160 (
            .O(N__31394),
            .I(N__31380));
    Span4Mux_s2_h I__7159 (
            .O(N__31391),
            .I(N__31375));
    LocalMux I__7158 (
            .O(N__31388),
            .I(N__31375));
    InMux I__7157 (
            .O(N__31387),
            .I(N__31371));
    InMux I__7156 (
            .O(N__31384),
            .I(N__31365));
    InMux I__7155 (
            .O(N__31383),
            .I(N__31361));
    Span4Mux_h I__7154 (
            .O(N__31380),
            .I(N__31356));
    Span4Mux_v I__7153 (
            .O(N__31375),
            .I(N__31356));
    InMux I__7152 (
            .O(N__31374),
            .I(N__31353));
    LocalMux I__7151 (
            .O(N__31371),
            .I(N__31348));
    InMux I__7150 (
            .O(N__31370),
            .I(N__31345));
    InMux I__7149 (
            .O(N__31369),
            .I(N__31342));
    InMux I__7148 (
            .O(N__31368),
            .I(N__31339));
    LocalMux I__7147 (
            .O(N__31365),
            .I(N__31336));
    InMux I__7146 (
            .O(N__31364),
            .I(N__31333));
    LocalMux I__7145 (
            .O(N__31361),
            .I(N__31325));
    Span4Mux_h I__7144 (
            .O(N__31356),
            .I(N__31325));
    LocalMux I__7143 (
            .O(N__31353),
            .I(N__31325));
    InMux I__7142 (
            .O(N__31352),
            .I(N__31319));
    InMux I__7141 (
            .O(N__31351),
            .I(N__31316));
    Span4Mux_v I__7140 (
            .O(N__31348),
            .I(N__31311));
    LocalMux I__7139 (
            .O(N__31345),
            .I(N__31311));
    LocalMux I__7138 (
            .O(N__31342),
            .I(N__31306));
    LocalMux I__7137 (
            .O(N__31339),
            .I(N__31306));
    Span4Mux_v I__7136 (
            .O(N__31336),
            .I(N__31303));
    LocalMux I__7135 (
            .O(N__31333),
            .I(N__31300));
    InMux I__7134 (
            .O(N__31332),
            .I(N__31297));
    Span4Mux_h I__7133 (
            .O(N__31325),
            .I(N__31294));
    CascadeMux I__7132 (
            .O(N__31324),
            .I(N__31291));
    InMux I__7131 (
            .O(N__31323),
            .I(N__31288));
    InMux I__7130 (
            .O(N__31322),
            .I(N__31285));
    LocalMux I__7129 (
            .O(N__31319),
            .I(N__31282));
    LocalMux I__7128 (
            .O(N__31316),
            .I(N__31275));
    Span4Mux_v I__7127 (
            .O(N__31311),
            .I(N__31275));
    Span4Mux_h I__7126 (
            .O(N__31306),
            .I(N__31275));
    Span4Mux_h I__7125 (
            .O(N__31303),
            .I(N__31270));
    Span4Mux_v I__7124 (
            .O(N__31300),
            .I(N__31270));
    LocalMux I__7123 (
            .O(N__31297),
            .I(N__31267));
    Span4Mux_s1_h I__7122 (
            .O(N__31294),
            .I(N__31264));
    InMux I__7121 (
            .O(N__31291),
            .I(N__31261));
    LocalMux I__7120 (
            .O(N__31288),
            .I(N__31258));
    LocalMux I__7119 (
            .O(N__31285),
            .I(N__31251));
    Span4Mux_h I__7118 (
            .O(N__31282),
            .I(N__31251));
    Span4Mux_h I__7117 (
            .O(N__31275),
            .I(N__31251));
    IoSpan4Mux I__7116 (
            .O(N__31270),
            .I(N__31248));
    Span4Mux_h I__7115 (
            .O(N__31267),
            .I(N__31243));
    Span4Mux_v I__7114 (
            .O(N__31264),
            .I(N__31243));
    LocalMux I__7113 (
            .O(N__31261),
            .I(cmd_13));
    Odrv12 I__7112 (
            .O(N__31258),
            .I(cmd_13));
    Odrv4 I__7111 (
            .O(N__31251),
            .I(cmd_13));
    Odrv4 I__7110 (
            .O(N__31248),
            .I(cmd_13));
    Odrv4 I__7109 (
            .O(N__31243),
            .I(cmd_13));
    InMux I__7108 (
            .O(N__31232),
            .I(N__31229));
    LocalMux I__7107 (
            .O(N__31229),
            .I(N__31226));
    Odrv4 I__7106 (
            .O(N__31226),
            .I(\Inst_core.Inst_sampler.n35 ));
    CascadeMux I__7105 (
            .O(N__31223),
            .I(N__31220));
    InMux I__7104 (
            .O(N__31220),
            .I(N__31217));
    LocalMux I__7103 (
            .O(N__31217),
            .I(N__31214));
    Odrv12 I__7102 (
            .O(N__31214),
            .I(\Inst_core.Inst_sampler.n36 ));
    InMux I__7101 (
            .O(N__31211),
            .I(N__31208));
    LocalMux I__7100 (
            .O(N__31208),
            .I(N__31205));
    Span4Mux_s2_h I__7099 (
            .O(N__31205),
            .I(N__31202));
    Odrv4 I__7098 (
            .O(N__31202),
            .I(\Inst_core.Inst_sampler.n33 ));
    CascadeMux I__7097 (
            .O(N__31199),
            .I(N__31193));
    InMux I__7096 (
            .O(N__31198),
            .I(N__31189));
    InMux I__7095 (
            .O(N__31197),
            .I(N__31186));
    InMux I__7094 (
            .O(N__31196),
            .I(N__31182));
    InMux I__7093 (
            .O(N__31193),
            .I(N__31177));
    InMux I__7092 (
            .O(N__31192),
            .I(N__31177));
    LocalMux I__7091 (
            .O(N__31189),
            .I(N__31172));
    LocalMux I__7090 (
            .O(N__31186),
            .I(N__31172));
    InMux I__7089 (
            .O(N__31185),
            .I(N__31169));
    LocalMux I__7088 (
            .O(N__31182),
            .I(N__31158));
    LocalMux I__7087 (
            .O(N__31177),
            .I(N__31158));
    Span4Mux_v I__7086 (
            .O(N__31172),
            .I(N__31153));
    LocalMux I__7085 (
            .O(N__31169),
            .I(N__31153));
    InMux I__7084 (
            .O(N__31168),
            .I(N__31146));
    InMux I__7083 (
            .O(N__31167),
            .I(N__31146));
    InMux I__7082 (
            .O(N__31166),
            .I(N__31146));
    InMux I__7081 (
            .O(N__31165),
            .I(N__31141));
    InMux I__7080 (
            .O(N__31164),
            .I(N__31141));
    InMux I__7079 (
            .O(N__31163),
            .I(N__31133));
    Span4Mux_v I__7078 (
            .O(N__31158),
            .I(N__31124));
    Span4Mux_h I__7077 (
            .O(N__31153),
            .I(N__31124));
    LocalMux I__7076 (
            .O(N__31146),
            .I(N__31124));
    LocalMux I__7075 (
            .O(N__31141),
            .I(N__31124));
    InMux I__7074 (
            .O(N__31140),
            .I(N__31115));
    InMux I__7073 (
            .O(N__31139),
            .I(N__31115));
    InMux I__7072 (
            .O(N__31138),
            .I(N__31115));
    InMux I__7071 (
            .O(N__31137),
            .I(N__31115));
    CascadeMux I__7070 (
            .O(N__31136),
            .I(N__31107));
    LocalMux I__7069 (
            .O(N__31133),
            .I(N__31099));
    Span4Mux_v I__7068 (
            .O(N__31124),
            .I(N__31094));
    LocalMux I__7067 (
            .O(N__31115),
            .I(N__31094));
    InMux I__7066 (
            .O(N__31114),
            .I(N__31082));
    InMux I__7065 (
            .O(N__31113),
            .I(N__31082));
    InMux I__7064 (
            .O(N__31112),
            .I(N__31082));
    InMux I__7063 (
            .O(N__31111),
            .I(N__31077));
    InMux I__7062 (
            .O(N__31110),
            .I(N__31077));
    InMux I__7061 (
            .O(N__31107),
            .I(N__31072));
    InMux I__7060 (
            .O(N__31106),
            .I(N__31072));
    InMux I__7059 (
            .O(N__31105),
            .I(N__31067));
    InMux I__7058 (
            .O(N__31104),
            .I(N__31067));
    InMux I__7057 (
            .O(N__31103),
            .I(N__31062));
    InMux I__7056 (
            .O(N__31102),
            .I(N__31062));
    Span4Mux_v I__7055 (
            .O(N__31099),
            .I(N__31057));
    Span4Mux_s3_v I__7054 (
            .O(N__31094),
            .I(N__31057));
    InMux I__7053 (
            .O(N__31093),
            .I(N__31054));
    InMux I__7052 (
            .O(N__31092),
            .I(N__31051));
    InMux I__7051 (
            .O(N__31091),
            .I(N__31048));
    InMux I__7050 (
            .O(N__31090),
            .I(N__31043));
    InMux I__7049 (
            .O(N__31089),
            .I(N__31043));
    LocalMux I__7048 (
            .O(N__31082),
            .I(N__31040));
    LocalMux I__7047 (
            .O(N__31077),
            .I(N__31035));
    LocalMux I__7046 (
            .O(N__31072),
            .I(N__31035));
    LocalMux I__7045 (
            .O(N__31067),
            .I(N__31032));
    LocalMux I__7044 (
            .O(N__31062),
            .I(N__31028));
    Span4Mux_h I__7043 (
            .O(N__31057),
            .I(N__31023));
    LocalMux I__7042 (
            .O(N__31054),
            .I(N__31023));
    LocalMux I__7041 (
            .O(N__31051),
            .I(N__31016));
    LocalMux I__7040 (
            .O(N__31048),
            .I(N__31016));
    LocalMux I__7039 (
            .O(N__31043),
            .I(N__31016));
    Span4Mux_v I__7038 (
            .O(N__31040),
            .I(N__31013));
    Span4Mux_v I__7037 (
            .O(N__31035),
            .I(N__31008));
    Span4Mux_v I__7036 (
            .O(N__31032),
            .I(N__31008));
    InMux I__7035 (
            .O(N__31031),
            .I(N__31005));
    Sp12to4 I__7034 (
            .O(N__31028),
            .I(N__30998));
    Sp12to4 I__7033 (
            .O(N__31023),
            .I(N__30998));
    Sp12to4 I__7032 (
            .O(N__31016),
            .I(N__30998));
    Span4Mux_h I__7031 (
            .O(N__31013),
            .I(N__30993));
    Span4Mux_v I__7030 (
            .O(N__31008),
            .I(N__30993));
    LocalMux I__7029 (
            .O(N__31005),
            .I(N__30987));
    Span12Mux_v I__7028 (
            .O(N__30998),
            .I(N__30987));
    Span4Mux_v I__7027 (
            .O(N__30993),
            .I(N__30984));
    InMux I__7026 (
            .O(N__30992),
            .I(N__30981));
    Odrv12 I__7025 (
            .O(N__30987),
            .I(wrDivider));
    Odrv4 I__7024 (
            .O(N__30984),
            .I(wrDivider));
    LocalMux I__7023 (
            .O(N__30981),
            .I(wrDivider));
    InMux I__7022 (
            .O(N__30974),
            .I(N__30971));
    LocalMux I__7021 (
            .O(N__30971),
            .I(N__30968));
    Span4Mux_s2_v I__7020 (
            .O(N__30968),
            .I(N__30965));
    Odrv4 I__7019 (
            .O(N__30965),
            .I(\Inst_core.Inst_sampler.n8669 ));
    CascadeMux I__7018 (
            .O(N__30962),
            .I(N__30959));
    InMux I__7017 (
            .O(N__30959),
            .I(N__30956));
    LocalMux I__7016 (
            .O(N__30956),
            .I(N__30953));
    Odrv4 I__7015 (
            .O(N__30953),
            .I(\Inst_core.Inst_sampler.n8671 ));
    InMux I__7014 (
            .O(N__30950),
            .I(N__30947));
    LocalMux I__7013 (
            .O(N__30947),
            .I(N__30944));
    Odrv4 I__7012 (
            .O(N__30944),
            .I(\Inst_core.Inst_sampler.n8673 ));
    CascadeMux I__7011 (
            .O(N__30941),
            .I(N__30937));
    InMux I__7010 (
            .O(N__30940),
            .I(N__30932));
    InMux I__7009 (
            .O(N__30937),
            .I(N__30929));
    InMux I__7008 (
            .O(N__30936),
            .I(N__30925));
    InMux I__7007 (
            .O(N__30935),
            .I(N__30918));
    LocalMux I__7006 (
            .O(N__30932),
            .I(N__30913));
    LocalMux I__7005 (
            .O(N__30929),
            .I(N__30913));
    InMux I__7004 (
            .O(N__30928),
            .I(N__30910));
    LocalMux I__7003 (
            .O(N__30925),
            .I(N__30906));
    InMux I__7002 (
            .O(N__30924),
            .I(N__30903));
    InMux I__7001 (
            .O(N__30923),
            .I(N__30900));
    InMux I__7000 (
            .O(N__30922),
            .I(N__30895));
    InMux I__6999 (
            .O(N__30921),
            .I(N__30895));
    LocalMux I__6998 (
            .O(N__30918),
            .I(N__30892));
    Span4Mux_v I__6997 (
            .O(N__30913),
            .I(N__30889));
    LocalMux I__6996 (
            .O(N__30910),
            .I(N__30886));
    InMux I__6995 (
            .O(N__30909),
            .I(N__30883));
    Span4Mux_v I__6994 (
            .O(N__30906),
            .I(N__30880));
    LocalMux I__6993 (
            .O(N__30903),
            .I(N__30875));
    LocalMux I__6992 (
            .O(N__30900),
            .I(N__30875));
    LocalMux I__6991 (
            .O(N__30895),
            .I(N__30872));
    Span4Mux_v I__6990 (
            .O(N__30892),
            .I(N__30867));
    Span4Mux_h I__6989 (
            .O(N__30889),
            .I(N__30867));
    Span12Mux_v I__6988 (
            .O(N__30886),
            .I(N__30864));
    LocalMux I__6987 (
            .O(N__30883),
            .I(N__30859));
    Span4Mux_v I__6986 (
            .O(N__30880),
            .I(N__30859));
    Span4Mux_v I__6985 (
            .O(N__30875),
            .I(N__30854));
    Span4Mux_h I__6984 (
            .O(N__30872),
            .I(N__30854));
    Odrv4 I__6983 (
            .O(N__30867),
            .I(memoryOut_2));
    Odrv12 I__6982 (
            .O(N__30864),
            .I(memoryOut_2));
    Odrv4 I__6981 (
            .O(N__30859),
            .I(memoryOut_2));
    Odrv4 I__6980 (
            .O(N__30854),
            .I(memoryOut_2));
    InMux I__6979 (
            .O(N__30845),
            .I(N__30842));
    LocalMux I__6978 (
            .O(N__30842),
            .I(N__30839));
    Span4Mux_s2_h I__6977 (
            .O(N__30839),
            .I(N__30835));
    InMux I__6976 (
            .O(N__30838),
            .I(N__30832));
    Odrv4 I__6975 (
            .O(N__30835),
            .I(valueRegister_2_adj_1334));
    LocalMux I__6974 (
            .O(N__30832),
            .I(valueRegister_2_adj_1334));
    InMux I__6973 (
            .O(N__30827),
            .I(N__30824));
    LocalMux I__6972 (
            .O(N__30824),
            .I(N__30820));
    CascadeMux I__6971 (
            .O(N__30823),
            .I(N__30817));
    Span4Mux_h I__6970 (
            .O(N__30820),
            .I(N__30813));
    InMux I__6969 (
            .O(N__30817),
            .I(N__30808));
    InMux I__6968 (
            .O(N__30816),
            .I(N__30808));
    Odrv4 I__6967 (
            .O(N__30813),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2 ));
    LocalMux I__6966 (
            .O(N__30808),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2 ));
    SRMux I__6965 (
            .O(N__30803),
            .I(N__30800));
    LocalMux I__6964 (
            .O(N__30800),
            .I(N__30797));
    Span4Mux_v I__6963 (
            .O(N__30797),
            .I(N__30794));
    Span4Mux_h I__6962 (
            .O(N__30794),
            .I(N__30791));
    Span4Mux_v I__6961 (
            .O(N__30791),
            .I(N__30788));
    Odrv4 I__6960 (
            .O(N__30788),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4754 ));
    InMux I__6959 (
            .O(N__30785),
            .I(N__30781));
    InMux I__6958 (
            .O(N__30784),
            .I(N__30778));
    LocalMux I__6957 (
            .O(N__30781),
            .I(N__30775));
    LocalMux I__6956 (
            .O(N__30778),
            .I(N__30772));
    Span4Mux_h I__6955 (
            .O(N__30775),
            .I(N__30768));
    Span4Mux_v I__6954 (
            .O(N__30772),
            .I(N__30765));
    InMux I__6953 (
            .O(N__30771),
            .I(N__30762));
    Span4Mux_v I__6952 (
            .O(N__30768),
            .I(N__30759));
    Span4Mux_h I__6951 (
            .O(N__30765),
            .I(N__30756));
    LocalMux I__6950 (
            .O(N__30762),
            .I(divider_11));
    Odrv4 I__6949 (
            .O(N__30759),
            .I(divider_11));
    Odrv4 I__6948 (
            .O(N__30756),
            .I(divider_11));
    InMux I__6947 (
            .O(N__30749),
            .I(N__30746));
    LocalMux I__6946 (
            .O(N__30746),
            .I(N__30742));
    InMux I__6945 (
            .O(N__30745),
            .I(N__30739));
    Span4Mux_s2_h I__6944 (
            .O(N__30742),
            .I(N__30736));
    LocalMux I__6943 (
            .O(N__30739),
            .I(\Inst_core.Inst_sampler.counter_23 ));
    Odrv4 I__6942 (
            .O(N__30736),
            .I(\Inst_core.Inst_sampler.counter_23 ));
    CascadeMux I__6941 (
            .O(N__30731),
            .I(N__30728));
    InMux I__6940 (
            .O(N__30728),
            .I(N__30722));
    InMux I__6939 (
            .O(N__30727),
            .I(N__30722));
    LocalMux I__6938 (
            .O(N__30722),
            .I(N__30718));
    InMux I__6937 (
            .O(N__30721),
            .I(N__30715));
    Span4Mux_v I__6936 (
            .O(N__30718),
            .I(N__30712));
    LocalMux I__6935 (
            .O(N__30715),
            .I(\Inst_core.Inst_sampler.counter_11 ));
    Odrv4 I__6934 (
            .O(N__30712),
            .I(\Inst_core.Inst_sampler.counter_11 ));
    InMux I__6933 (
            .O(N__30707),
            .I(N__30704));
    LocalMux I__6932 (
            .O(N__30704),
            .I(N__30700));
    InMux I__6931 (
            .O(N__30703),
            .I(N__30696));
    Span4Mux_s2_h I__6930 (
            .O(N__30700),
            .I(N__30693));
    InMux I__6929 (
            .O(N__30699),
            .I(N__30690));
    LocalMux I__6928 (
            .O(N__30696),
            .I(\Inst_core.Inst_sampler.counter_2 ));
    Odrv4 I__6927 (
            .O(N__30693),
            .I(\Inst_core.Inst_sampler.counter_2 ));
    LocalMux I__6926 (
            .O(N__30690),
            .I(\Inst_core.Inst_sampler.counter_2 ));
    InMux I__6925 (
            .O(N__30683),
            .I(N__30680));
    LocalMux I__6924 (
            .O(N__30680),
            .I(N__30677));
    Odrv4 I__6923 (
            .O(N__30677),
            .I(\Inst_core.Inst_sampler.n8606 ));
    CascadeMux I__6922 (
            .O(N__30674),
            .I(\Inst_core.Inst_sampler.n3_cascade_ ));
    CascadeMux I__6921 (
            .O(N__30671),
            .I(N__30667));
    InMux I__6920 (
            .O(N__30670),
            .I(N__30661));
    InMux I__6919 (
            .O(N__30667),
            .I(N__30661));
    InMux I__6918 (
            .O(N__30666),
            .I(N__30658));
    LocalMux I__6917 (
            .O(N__30661),
            .I(N__30655));
    LocalMux I__6916 (
            .O(N__30658),
            .I(divider_23));
    Odrv12 I__6915 (
            .O(N__30655),
            .I(divider_23));
    InMux I__6914 (
            .O(N__30650),
            .I(N__30647));
    LocalMux I__6913 (
            .O(N__30647),
            .I(N__30644));
    Odrv4 I__6912 (
            .O(N__30644),
            .I(\Inst_core.Inst_sampler.n8618 ));
    CascadeMux I__6911 (
            .O(N__30641),
            .I(\Inst_core.Inst_sampler.n8656_cascade_ ));
    InMux I__6910 (
            .O(N__30638),
            .I(N__30633));
    InMux I__6909 (
            .O(N__30637),
            .I(N__30630));
    InMux I__6908 (
            .O(N__30636),
            .I(N__30627));
    LocalMux I__6907 (
            .O(N__30633),
            .I(N__30622));
    LocalMux I__6906 (
            .O(N__30630),
            .I(N__30622));
    LocalMux I__6905 (
            .O(N__30627),
            .I(divider_1));
    Odrv12 I__6904 (
            .O(N__30622),
            .I(divider_1));
    InMux I__6903 (
            .O(N__30617),
            .I(N__30613));
    InMux I__6902 (
            .O(N__30616),
            .I(N__30610));
    LocalMux I__6901 (
            .O(N__30613),
            .I(N__30606));
    LocalMux I__6900 (
            .O(N__30610),
            .I(N__30603));
    InMux I__6899 (
            .O(N__30609),
            .I(N__30600));
    Span4Mux_v I__6898 (
            .O(N__30606),
            .I(N__30595));
    Span4Mux_v I__6897 (
            .O(N__30603),
            .I(N__30595));
    LocalMux I__6896 (
            .O(N__30600),
            .I(\Inst_core.Inst_sampler.counter_18 ));
    Odrv4 I__6895 (
            .O(N__30595),
            .I(\Inst_core.Inst_sampler.counter_18 ));
    CascadeMux I__6894 (
            .O(N__30590),
            .I(N__30587));
    InMux I__6893 (
            .O(N__30587),
            .I(N__30584));
    LocalMux I__6892 (
            .O(N__30584),
            .I(N__30580));
    InMux I__6891 (
            .O(N__30583),
            .I(N__30576));
    Span4Mux_v I__6890 (
            .O(N__30580),
            .I(N__30573));
    InMux I__6889 (
            .O(N__30579),
            .I(N__30570));
    LocalMux I__6888 (
            .O(N__30576),
            .I(N__30567));
    Span4Mux_s0_h I__6887 (
            .O(N__30573),
            .I(N__30564));
    LocalMux I__6886 (
            .O(N__30570),
            .I(divider_18));
    Odrv4 I__6885 (
            .O(N__30567),
            .I(divider_18));
    Odrv4 I__6884 (
            .O(N__30564),
            .I(divider_18));
    InMux I__6883 (
            .O(N__30557),
            .I(N__30552));
    InMux I__6882 (
            .O(N__30556),
            .I(N__30549));
    InMux I__6881 (
            .O(N__30555),
            .I(N__30546));
    LocalMux I__6880 (
            .O(N__30552),
            .I(N__30541));
    LocalMux I__6879 (
            .O(N__30549),
            .I(N__30541));
    LocalMux I__6878 (
            .O(N__30546),
            .I(\Inst_core.Inst_sampler.counter_1 ));
    Odrv4 I__6877 (
            .O(N__30541),
            .I(\Inst_core.Inst_sampler.counter_1 ));
    InMux I__6876 (
            .O(N__30536),
            .I(N__30533));
    LocalMux I__6875 (
            .O(N__30533),
            .I(N__30530));
    Odrv4 I__6874 (
            .O(N__30530),
            .I(\Inst_core.Inst_sampler.n28 ));
    CascadeMux I__6873 (
            .O(N__30527),
            .I(\Inst_core.Inst_sampler.n27_cascade_ ));
    InMux I__6872 (
            .O(N__30524),
            .I(N__30519));
    InMux I__6871 (
            .O(N__30523),
            .I(N__30516));
    InMux I__6870 (
            .O(N__30522),
            .I(N__30513));
    LocalMux I__6869 (
            .O(N__30519),
            .I(N__30508));
    LocalMux I__6868 (
            .O(N__30516),
            .I(N__30508));
    LocalMux I__6867 (
            .O(N__30513),
            .I(divider_6));
    Odrv12 I__6866 (
            .O(N__30508),
            .I(divider_6));
    InMux I__6865 (
            .O(N__30503),
            .I(N__30498));
    InMux I__6864 (
            .O(N__30502),
            .I(N__30495));
    InMux I__6863 (
            .O(N__30501),
            .I(N__30492));
    LocalMux I__6862 (
            .O(N__30498),
            .I(N__30487));
    LocalMux I__6861 (
            .O(N__30495),
            .I(N__30487));
    LocalMux I__6860 (
            .O(N__30492),
            .I(\Inst_core.Inst_sampler.counter_3 ));
    Odrv4 I__6859 (
            .O(N__30487),
            .I(\Inst_core.Inst_sampler.counter_3 ));
    SRMux I__6858 (
            .O(N__30482),
            .I(N__30479));
    LocalMux I__6857 (
            .O(N__30479),
            .I(N__30476));
    Span4Mux_v I__6856 (
            .O(N__30476),
            .I(N__30473));
    Span4Mux_h I__6855 (
            .O(N__30473),
            .I(N__30470));
    Odrv4 I__6854 (
            .O(N__30470),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4747 ));
    CascadeMux I__6853 (
            .O(N__30467),
            .I(N__30463));
    CascadeMux I__6852 (
            .O(N__30466),
            .I(N__30458));
    InMux I__6851 (
            .O(N__30463),
            .I(N__30453));
    InMux I__6850 (
            .O(N__30462),
            .I(N__30449));
    InMux I__6849 (
            .O(N__30461),
            .I(N__30446));
    InMux I__6848 (
            .O(N__30458),
            .I(N__30443));
    InMux I__6847 (
            .O(N__30457),
            .I(N__30439));
    InMux I__6846 (
            .O(N__30456),
            .I(N__30436));
    LocalMux I__6845 (
            .O(N__30453),
            .I(N__30433));
    InMux I__6844 (
            .O(N__30452),
            .I(N__30429));
    LocalMux I__6843 (
            .O(N__30449),
            .I(N__30426));
    LocalMux I__6842 (
            .O(N__30446),
            .I(N__30423));
    LocalMux I__6841 (
            .O(N__30443),
            .I(N__30420));
    InMux I__6840 (
            .O(N__30442),
            .I(N__30417));
    LocalMux I__6839 (
            .O(N__30439),
            .I(N__30414));
    LocalMux I__6838 (
            .O(N__30436),
            .I(N__30409));
    Span4Mux_h I__6837 (
            .O(N__30433),
            .I(N__30409));
    InMux I__6836 (
            .O(N__30432),
            .I(N__30406));
    LocalMux I__6835 (
            .O(N__30429),
            .I(N__30402));
    Span4Mux_v I__6834 (
            .O(N__30426),
            .I(N__30397));
    Span4Mux_s3_v I__6833 (
            .O(N__30423),
            .I(N__30397));
    Span4Mux_h I__6832 (
            .O(N__30420),
            .I(N__30394));
    LocalMux I__6831 (
            .O(N__30417),
            .I(N__30391));
    Sp12to4 I__6830 (
            .O(N__30414),
            .I(N__30386));
    Sp12to4 I__6829 (
            .O(N__30409),
            .I(N__30386));
    LocalMux I__6828 (
            .O(N__30406),
            .I(N__30383));
    InMux I__6827 (
            .O(N__30405),
            .I(N__30380));
    Span4Mux_h I__6826 (
            .O(N__30402),
            .I(N__30373));
    Span4Mux_h I__6825 (
            .O(N__30397),
            .I(N__30373));
    Span4Mux_v I__6824 (
            .O(N__30394),
            .I(N__30373));
    Span12Mux_s5_h I__6823 (
            .O(N__30391),
            .I(N__30366));
    Span12Mux_s11_v I__6822 (
            .O(N__30386),
            .I(N__30366));
    Span12Mux_s6_h I__6821 (
            .O(N__30383),
            .I(N__30366));
    LocalMux I__6820 (
            .O(N__30380),
            .I(memoryOut_6));
    Odrv4 I__6819 (
            .O(N__30373),
            .I(memoryOut_6));
    Odrv12 I__6818 (
            .O(N__30366),
            .I(memoryOut_6));
    InMux I__6817 (
            .O(N__30359),
            .I(N__30354));
    InMux I__6816 (
            .O(N__30358),
            .I(N__30351));
    CascadeMux I__6815 (
            .O(N__30357),
            .I(N__30348));
    LocalMux I__6814 (
            .O(N__30354),
            .I(N__30339));
    LocalMux I__6813 (
            .O(N__30351),
            .I(N__30339));
    InMux I__6812 (
            .O(N__30348),
            .I(N__30336));
    CascadeMux I__6811 (
            .O(N__30347),
            .I(N__30333));
    CascadeMux I__6810 (
            .O(N__30346),
            .I(N__30329));
    InMux I__6809 (
            .O(N__30345),
            .I(N__30326));
    InMux I__6808 (
            .O(N__30344),
            .I(N__30323));
    Span4Mux_h I__6807 (
            .O(N__30339),
            .I(N__30320));
    LocalMux I__6806 (
            .O(N__30336),
            .I(N__30317));
    InMux I__6805 (
            .O(N__30333),
            .I(N__30314));
    InMux I__6804 (
            .O(N__30332),
            .I(N__30311));
    InMux I__6803 (
            .O(N__30329),
            .I(N__30308));
    LocalMux I__6802 (
            .O(N__30326),
            .I(N__30305));
    LocalMux I__6801 (
            .O(N__30323),
            .I(N__30302));
    Span4Mux_h I__6800 (
            .O(N__30320),
            .I(N__30297));
    Span4Mux_h I__6799 (
            .O(N__30317),
            .I(N__30297));
    LocalMux I__6798 (
            .O(N__30314),
            .I(N__30293));
    LocalMux I__6797 (
            .O(N__30311),
            .I(N__30288));
    LocalMux I__6796 (
            .O(N__30308),
            .I(N__30288));
    Span4Mux_s2_v I__6795 (
            .O(N__30305),
            .I(N__30285));
    Span4Mux_s2_h I__6794 (
            .O(N__30302),
            .I(N__30282));
    Span4Mux_v I__6793 (
            .O(N__30297),
            .I(N__30279));
    InMux I__6792 (
            .O(N__30296),
            .I(N__30276));
    Span4Mux_v I__6791 (
            .O(N__30293),
            .I(N__30273));
    Span4Mux_v I__6790 (
            .O(N__30288),
            .I(N__30268));
    Span4Mux_v I__6789 (
            .O(N__30285),
            .I(N__30268));
    Span4Mux_v I__6788 (
            .O(N__30282),
            .I(N__30263));
    Span4Mux_h I__6787 (
            .O(N__30279),
            .I(N__30263));
    LocalMux I__6786 (
            .O(N__30276),
            .I(configRegister_26_adj_1297));
    Odrv4 I__6785 (
            .O(N__30273),
            .I(configRegister_26_adj_1297));
    Odrv4 I__6784 (
            .O(N__30268),
            .I(configRegister_26_adj_1297));
    Odrv4 I__6783 (
            .O(N__30263),
            .I(configRegister_26_adj_1297));
    InMux I__6782 (
            .O(N__30254),
            .I(N__30251));
    LocalMux I__6781 (
            .O(N__30251),
            .I(N__30248));
    Span4Mux_s2_h I__6780 (
            .O(N__30248),
            .I(N__30245));
    Span4Mux_h I__6779 (
            .O(N__30245),
            .I(N__30241));
    InMux I__6778 (
            .O(N__30244),
            .I(N__30238));
    Odrv4 I__6777 (
            .O(N__30241),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6 ));
    LocalMux I__6776 (
            .O(N__30238),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6 ));
    InMux I__6775 (
            .O(N__30233),
            .I(N__30230));
    LocalMux I__6774 (
            .O(N__30230),
            .I(N__30227));
    Span4Mux_v I__6773 (
            .O(N__30227),
            .I(N__30224));
    Odrv4 I__6772 (
            .O(N__30224),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_6 ));
    SRMux I__6771 (
            .O(N__30221),
            .I(N__30218));
    LocalMux I__6770 (
            .O(N__30218),
            .I(N__30215));
    Span4Mux_v I__6769 (
            .O(N__30215),
            .I(N__30212));
    Odrv4 I__6768 (
            .O(N__30212),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4751 ));
    InMux I__6767 (
            .O(N__30209),
            .I(N__30206));
    LocalMux I__6766 (
            .O(N__30206),
            .I(N__30202));
    InMux I__6765 (
            .O(N__30205),
            .I(N__30199));
    Span4Mux_v I__6764 (
            .O(N__30202),
            .I(N__30196));
    LocalMux I__6763 (
            .O(N__30199),
            .I(fwd_0));
    Odrv4 I__6762 (
            .O(N__30196),
            .I(fwd_0));
    CascadeMux I__6761 (
            .O(N__30191),
            .I(N__30188));
    InMux I__6760 (
            .O(N__30188),
            .I(N__30184));
    InMux I__6759 (
            .O(N__30187),
            .I(N__30181));
    LocalMux I__6758 (
            .O(N__30184),
            .I(N__30178));
    LocalMux I__6757 (
            .O(N__30181),
            .I(fwd_2));
    Odrv12 I__6756 (
            .O(N__30178),
            .I(fwd_2));
    CascadeMux I__6755 (
            .O(N__30173),
            .I(N__30170));
    InMux I__6754 (
            .O(N__30170),
            .I(N__30167));
    LocalMux I__6753 (
            .O(N__30167),
            .I(N__30164));
    Span4Mux_v I__6752 (
            .O(N__30164),
            .I(N__30161));
    Span4Mux_h I__6751 (
            .O(N__30161),
            .I(N__30158));
    Odrv4 I__6750 (
            .O(N__30158),
            .I(\Inst_core.Inst_controller.n16 ));
    IoInMux I__6749 (
            .O(N__30155),
            .I(N__30151));
    InMux I__6748 (
            .O(N__30154),
            .I(N__30148));
    LocalMux I__6747 (
            .O(N__30151),
            .I(N__30145));
    LocalMux I__6746 (
            .O(N__30148),
            .I(N__30141));
    Span4Mux_s1_h I__6745 (
            .O(N__30145),
            .I(N__30138));
    InMux I__6744 (
            .O(N__30144),
            .I(N__30135));
    Span12Mux_s10_h I__6743 (
            .O(N__30141),
            .I(N__30132));
    Odrv4 I__6742 (
            .O(N__30138),
            .I(debugleds_c_1));
    LocalMux I__6741 (
            .O(N__30135),
            .I(debugleds_c_1));
    Odrv12 I__6740 (
            .O(N__30132),
            .I(debugleds_c_1));
    CascadeMux I__6739 (
            .O(N__30125),
            .I(\Inst_core.n4_cascade_ ));
    CascadeMux I__6738 (
            .O(N__30122),
            .I(\Inst_core.Inst_controller.n3907_cascade_ ));
    CascadeMux I__6737 (
            .O(N__30119),
            .I(N__30116));
    InMux I__6736 (
            .O(N__30116),
            .I(N__30110));
    InMux I__6735 (
            .O(N__30115),
            .I(N__30107));
    InMux I__6734 (
            .O(N__30114),
            .I(N__30104));
    CascadeMux I__6733 (
            .O(N__30113),
            .I(N__30101));
    LocalMux I__6732 (
            .O(N__30110),
            .I(N__30095));
    LocalMux I__6731 (
            .O(N__30107),
            .I(N__30095));
    LocalMux I__6730 (
            .O(N__30104),
            .I(N__30092));
    InMux I__6729 (
            .O(N__30101),
            .I(N__30089));
    InMux I__6728 (
            .O(N__30100),
            .I(N__30086));
    Span4Mux_h I__6727 (
            .O(N__30095),
            .I(N__30082));
    Span4Mux_h I__6726 (
            .O(N__30092),
            .I(N__30079));
    LocalMux I__6725 (
            .O(N__30089),
            .I(N__30076));
    LocalMux I__6724 (
            .O(N__30086),
            .I(N__30073));
    InMux I__6723 (
            .O(N__30085),
            .I(N__30070));
    Span4Mux_v I__6722 (
            .O(N__30082),
            .I(N__30065));
    Span4Mux_v I__6721 (
            .O(N__30079),
            .I(N__30062));
    Span4Mux_v I__6720 (
            .O(N__30076),
            .I(N__30059));
    Span4Mux_h I__6719 (
            .O(N__30073),
            .I(N__30054));
    LocalMux I__6718 (
            .O(N__30070),
            .I(N__30054));
    InMux I__6717 (
            .O(N__30069),
            .I(N__30051));
    InMux I__6716 (
            .O(N__30068),
            .I(N__30048));
    Odrv4 I__6715 (
            .O(N__30065),
            .I(cmd_22));
    Odrv4 I__6714 (
            .O(N__30062),
            .I(cmd_22));
    Odrv4 I__6713 (
            .O(N__30059),
            .I(cmd_22));
    Odrv4 I__6712 (
            .O(N__30054),
            .I(cmd_22));
    LocalMux I__6711 (
            .O(N__30051),
            .I(cmd_22));
    LocalMux I__6710 (
            .O(N__30048),
            .I(cmd_22));
    InMux I__6709 (
            .O(N__30035),
            .I(N__30030));
    CascadeMux I__6708 (
            .O(N__30034),
            .I(N__30027));
    CascadeMux I__6707 (
            .O(N__30033),
            .I(N__30024));
    LocalMux I__6706 (
            .O(N__30030),
            .I(N__30020));
    InMux I__6705 (
            .O(N__30027),
            .I(N__30017));
    InMux I__6704 (
            .O(N__30024),
            .I(N__30012));
    InMux I__6703 (
            .O(N__30023),
            .I(N__30012));
    Span4Mux_v I__6702 (
            .O(N__30020),
            .I(N__30009));
    LocalMux I__6701 (
            .O(N__30017),
            .I(cmd_26));
    LocalMux I__6700 (
            .O(N__30012),
            .I(cmd_26));
    Odrv4 I__6699 (
            .O(N__30009),
            .I(cmd_26));
    CascadeMux I__6698 (
            .O(N__30002),
            .I(N__29998));
    InMux I__6697 (
            .O(N__30001),
            .I(N__29993));
    InMux I__6696 (
            .O(N__29998),
            .I(N__29993));
    LocalMux I__6695 (
            .O(N__29993),
            .I(N__29990));
    Span4Mux_s2_h I__6694 (
            .O(N__29990),
            .I(N__29985));
    InMux I__6693 (
            .O(N__29989),
            .I(N__29980));
    InMux I__6692 (
            .O(N__29988),
            .I(N__29980));
    Odrv4 I__6691 (
            .O(N__29985),
            .I(cmd_27));
    LocalMux I__6690 (
            .O(N__29980),
            .I(cmd_27));
    CascadeMux I__6689 (
            .O(N__29975),
            .I(N__29972));
    InMux I__6688 (
            .O(N__29972),
            .I(N__29968));
    CascadeMux I__6687 (
            .O(N__29971),
            .I(N__29965));
    LocalMux I__6686 (
            .O(N__29968),
            .I(N__29962));
    InMux I__6685 (
            .O(N__29965),
            .I(N__29959));
    Span4Mux_h I__6684 (
            .O(N__29962),
            .I(N__29955));
    LocalMux I__6683 (
            .O(N__29959),
            .I(N__29952));
    InMux I__6682 (
            .O(N__29958),
            .I(N__29949));
    Span4Mux_v I__6681 (
            .O(N__29955),
            .I(N__29946));
    Span4Mux_h I__6680 (
            .O(N__29952),
            .I(N__29943));
    LocalMux I__6679 (
            .O(N__29949),
            .I(divider_19));
    Odrv4 I__6678 (
            .O(N__29946),
            .I(divider_19));
    Odrv4 I__6677 (
            .O(N__29943),
            .I(divider_19));
    InMux I__6676 (
            .O(N__29936),
            .I(N__29933));
    LocalMux I__6675 (
            .O(N__29933),
            .I(N__29929));
    InMux I__6674 (
            .O(N__29932),
            .I(N__29926));
    Span4Mux_s3_h I__6673 (
            .O(N__29929),
            .I(N__29923));
    LocalMux I__6672 (
            .O(N__29926),
            .I(bwd_2));
    Odrv4 I__6671 (
            .O(N__29923),
            .I(bwd_2));
    CascadeMux I__6670 (
            .O(N__29918),
            .I(N__29915));
    InMux I__6669 (
            .O(N__29915),
            .I(N__29911));
    InMux I__6668 (
            .O(N__29914),
            .I(N__29908));
    LocalMux I__6667 (
            .O(N__29911),
            .I(N__29905));
    LocalMux I__6666 (
            .O(N__29908),
            .I(bwd_13));
    Odrv12 I__6665 (
            .O(N__29905),
            .I(bwd_13));
    InMux I__6664 (
            .O(N__29900),
            .I(N__29897));
    LocalMux I__6663 (
            .O(N__29897),
            .I(N__29894));
    Span4Mux_s3_h I__6662 (
            .O(N__29894),
            .I(N__29891));
    Odrv4 I__6661 (
            .O(N__29891),
            .I(\Inst_core.Inst_controller.n18_adj_990 ));
    InMux I__6660 (
            .O(N__29888),
            .I(N__29885));
    LocalMux I__6659 (
            .O(N__29885),
            .I(N__29882));
    Odrv12 I__6658 (
            .O(N__29882),
            .I(\Inst_core.Inst_controller.n20 ));
    CascadeMux I__6657 (
            .O(N__29879),
            .I(\Inst_core.Inst_controller.n17_cascade_ ));
    InMux I__6656 (
            .O(N__29876),
            .I(N__29873));
    LocalMux I__6655 (
            .O(N__29873),
            .I(N__29870));
    Span4Mux_s2_h I__6654 (
            .O(N__29870),
            .I(N__29867));
    Odrv4 I__6653 (
            .O(N__29867),
            .I(\Inst_core.Inst_controller.n30 ));
    CascadeMux I__6652 (
            .O(N__29864),
            .I(\Inst_core.Inst_controller.n29_cascade_ ));
    InMux I__6651 (
            .O(N__29861),
            .I(N__29858));
    LocalMux I__6650 (
            .O(N__29858),
            .I(N__29855));
    Span4Mux_h I__6649 (
            .O(N__29855),
            .I(N__29852));
    Odrv4 I__6648 (
            .O(N__29852),
            .I(\Inst_core.Inst_controller.n6693 ));
    InMux I__6647 (
            .O(N__29849),
            .I(N__29845));
    InMux I__6646 (
            .O(N__29848),
            .I(N__29842));
    LocalMux I__6645 (
            .O(N__29845),
            .I(N__29839));
    LocalMux I__6644 (
            .O(N__29842),
            .I(\Inst_core.Inst_controller.bwd_14 ));
    Odrv4 I__6643 (
            .O(N__29839),
            .I(\Inst_core.Inst_controller.bwd_14 ));
    InMux I__6642 (
            .O(N__29834),
            .I(N__29831));
    LocalMux I__6641 (
            .O(N__29831),
            .I(\Inst_core.Inst_controller.n19 ));
    InMux I__6640 (
            .O(N__29828),
            .I(N__29825));
    LocalMux I__6639 (
            .O(N__29825),
            .I(N__29821));
    InMux I__6638 (
            .O(N__29824),
            .I(N__29818));
    Odrv4 I__6637 (
            .O(N__29821),
            .I(valueRegister_2_adj_1294));
    LocalMux I__6636 (
            .O(N__29818),
            .I(valueRegister_2_adj_1294));
    InMux I__6635 (
            .O(N__29813),
            .I(N__29810));
    LocalMux I__6634 (
            .O(N__29810),
            .I(N__29806));
    CascadeMux I__6633 (
            .O(N__29809),
            .I(N__29803));
    Span4Mux_s2_h I__6632 (
            .O(N__29806),
            .I(N__29799));
    InMux I__6631 (
            .O(N__29803),
            .I(N__29794));
    InMux I__6630 (
            .O(N__29802),
            .I(N__29794));
    Odrv4 I__6629 (
            .O(N__29799),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2 ));
    LocalMux I__6628 (
            .O(N__29794),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2 ));
    InMux I__6627 (
            .O(N__29789),
            .I(N__29786));
    LocalMux I__6626 (
            .O(N__29786),
            .I(N__29783));
    Odrv12 I__6625 (
            .O(N__29783),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_2 ));
    InMux I__6624 (
            .O(N__29780),
            .I(N__29776));
    InMux I__6623 (
            .O(N__29779),
            .I(N__29773));
    LocalMux I__6622 (
            .O(N__29776),
            .I(N__29770));
    LocalMux I__6621 (
            .O(N__29773),
            .I(maskRegister_6_adj_1282));
    Odrv12 I__6620 (
            .O(N__29770),
            .I(maskRegister_6_adj_1282));
    InMux I__6619 (
            .O(N__29765),
            .I(N__29759));
    InMux I__6618 (
            .O(N__29764),
            .I(N__29759));
    LocalMux I__6617 (
            .O(N__29759),
            .I(N__29753));
    InMux I__6616 (
            .O(N__29758),
            .I(N__29746));
    InMux I__6615 (
            .O(N__29757),
            .I(N__29746));
    CascadeMux I__6614 (
            .O(N__29756),
            .I(N__29742));
    Span4Mux_v I__6613 (
            .O(N__29753),
            .I(N__29739));
    InMux I__6612 (
            .O(N__29752),
            .I(N__29736));
    InMux I__6611 (
            .O(N__29751),
            .I(N__29733));
    LocalMux I__6610 (
            .O(N__29746),
            .I(N__29730));
    InMux I__6609 (
            .O(N__29745),
            .I(N__29725));
    InMux I__6608 (
            .O(N__29742),
            .I(N__29725));
    Odrv4 I__6607 (
            .O(N__29739),
            .I(cmd_31));
    LocalMux I__6606 (
            .O(N__29736),
            .I(cmd_31));
    LocalMux I__6605 (
            .O(N__29733),
            .I(cmd_31));
    Odrv4 I__6604 (
            .O(N__29730),
            .I(cmd_31));
    LocalMux I__6603 (
            .O(N__29725),
            .I(cmd_31));
    InMux I__6602 (
            .O(N__29714),
            .I(N__29708));
    InMux I__6601 (
            .O(N__29713),
            .I(N__29699));
    InMux I__6600 (
            .O(N__29712),
            .I(N__29699));
    InMux I__6599 (
            .O(N__29711),
            .I(N__29699));
    LocalMux I__6598 (
            .O(N__29708),
            .I(N__29696));
    InMux I__6597 (
            .O(N__29707),
            .I(N__29693));
    InMux I__6596 (
            .O(N__29706),
            .I(N__29688));
    LocalMux I__6595 (
            .O(N__29699),
            .I(N__29685));
    Span4Mux_h I__6594 (
            .O(N__29696),
            .I(N__29680));
    LocalMux I__6593 (
            .O(N__29693),
            .I(N__29680));
    InMux I__6592 (
            .O(N__29692),
            .I(N__29672));
    CascadeMux I__6591 (
            .O(N__29691),
            .I(N__29668));
    LocalMux I__6590 (
            .O(N__29688),
            .I(N__29665));
    Span4Mux_v I__6589 (
            .O(N__29685),
            .I(N__29662));
    Span4Mux_v I__6588 (
            .O(N__29680),
            .I(N__29659));
    InMux I__6587 (
            .O(N__29679),
            .I(N__29656));
    InMux I__6586 (
            .O(N__29678),
            .I(N__29653));
    InMux I__6585 (
            .O(N__29677),
            .I(N__29650));
    InMux I__6584 (
            .O(N__29676),
            .I(N__29647));
    InMux I__6583 (
            .O(N__29675),
            .I(N__29644));
    LocalMux I__6582 (
            .O(N__29672),
            .I(N__29641));
    InMux I__6581 (
            .O(N__29671),
            .I(N__29638));
    InMux I__6580 (
            .O(N__29668),
            .I(N__29635));
    Span4Mux_v I__6579 (
            .O(N__29665),
            .I(N__29626));
    Span4Mux_h I__6578 (
            .O(N__29662),
            .I(N__29626));
    Span4Mux_s2_v I__6577 (
            .O(N__29659),
            .I(N__29626));
    LocalMux I__6576 (
            .O(N__29656),
            .I(N__29626));
    LocalMux I__6575 (
            .O(N__29653),
            .I(N__29616));
    LocalMux I__6574 (
            .O(N__29650),
            .I(N__29616));
    LocalMux I__6573 (
            .O(N__29647),
            .I(N__29616));
    LocalMux I__6572 (
            .O(N__29644),
            .I(N__29611));
    Span4Mux_v I__6571 (
            .O(N__29641),
            .I(N__29611));
    LocalMux I__6570 (
            .O(N__29638),
            .I(N__29606));
    LocalMux I__6569 (
            .O(N__29635),
            .I(N__29606));
    Sp12to4 I__6568 (
            .O(N__29626),
            .I(N__29603));
    InMux I__6567 (
            .O(N__29625),
            .I(N__29598));
    InMux I__6566 (
            .O(N__29624),
            .I(N__29598));
    InMux I__6565 (
            .O(N__29623),
            .I(N__29595));
    Span4Mux_v I__6564 (
            .O(N__29616),
            .I(N__29592));
    Span4Mux_h I__6563 (
            .O(N__29611),
            .I(N__29589));
    Span12Mux_s6_h I__6562 (
            .O(N__29606),
            .I(N__29584));
    Span12Mux_s7_v I__6561 (
            .O(N__29603),
            .I(N__29584));
    LocalMux I__6560 (
            .O(N__29598),
            .I(cmd_10));
    LocalMux I__6559 (
            .O(N__29595),
            .I(cmd_10));
    Odrv4 I__6558 (
            .O(N__29592),
            .I(cmd_10));
    Odrv4 I__6557 (
            .O(N__29589),
            .I(cmd_10));
    Odrv12 I__6556 (
            .O(N__29584),
            .I(cmd_10));
    CascadeMux I__6555 (
            .O(N__29573),
            .I(N__29570));
    InMux I__6554 (
            .O(N__29570),
            .I(N__29567));
    LocalMux I__6553 (
            .O(N__29567),
            .I(N__29563));
    InMux I__6552 (
            .O(N__29566),
            .I(N__29560));
    Odrv12 I__6551 (
            .O(N__29563),
            .I(valueRegister_2_adj_1374));
    LocalMux I__6550 (
            .O(N__29560),
            .I(valueRegister_2_adj_1374));
    InMux I__6549 (
            .O(N__29555),
            .I(N__29549));
    InMux I__6548 (
            .O(N__29554),
            .I(N__29549));
    LocalMux I__6547 (
            .O(N__29549),
            .I(N__29545));
    InMux I__6546 (
            .O(N__29548),
            .I(N__29542));
    Span4Mux_h I__6545 (
            .O(N__29545),
            .I(N__29535));
    LocalMux I__6544 (
            .O(N__29542),
            .I(N__29535));
    InMux I__6543 (
            .O(N__29541),
            .I(N__29532));
    InMux I__6542 (
            .O(N__29540),
            .I(N__29529));
    Span4Mux_s3_h I__6541 (
            .O(N__29535),
            .I(N__29520));
    LocalMux I__6540 (
            .O(N__29532),
            .I(N__29520));
    LocalMux I__6539 (
            .O(N__29529),
            .I(N__29520));
    InMux I__6538 (
            .O(N__29528),
            .I(N__29517));
    CascadeMux I__6537 (
            .O(N__29527),
            .I(N__29514));
    Span4Mux_v I__6536 (
            .O(N__29520),
            .I(N__29510));
    LocalMux I__6535 (
            .O(N__29517),
            .I(N__29507));
    InMux I__6534 (
            .O(N__29514),
            .I(N__29502));
    InMux I__6533 (
            .O(N__29513),
            .I(N__29502));
    Odrv4 I__6532 (
            .O(N__29510),
            .I(cmd_25));
    Odrv12 I__6531 (
            .O(N__29507),
            .I(cmd_25));
    LocalMux I__6530 (
            .O(N__29502),
            .I(cmd_25));
    CascadeMux I__6529 (
            .O(N__29495),
            .I(N__29491));
    InMux I__6528 (
            .O(N__29494),
            .I(N__29484));
    InMux I__6527 (
            .O(N__29491),
            .I(N__29484));
    InMux I__6526 (
            .O(N__29490),
            .I(N__29479));
    InMux I__6525 (
            .O(N__29489),
            .I(N__29476));
    LocalMux I__6524 (
            .O(N__29484),
            .I(N__29472));
    InMux I__6523 (
            .O(N__29483),
            .I(N__29467));
    InMux I__6522 (
            .O(N__29482),
            .I(N__29467));
    LocalMux I__6521 (
            .O(N__29479),
            .I(N__29464));
    LocalMux I__6520 (
            .O(N__29476),
            .I(N__29461));
    InMux I__6519 (
            .O(N__29475),
            .I(N__29458));
    Span4Mux_h I__6518 (
            .O(N__29472),
            .I(N__29452));
    LocalMux I__6517 (
            .O(N__29467),
            .I(N__29452));
    Span4Mux_v I__6516 (
            .O(N__29464),
            .I(N__29449));
    Span4Mux_s2_h I__6515 (
            .O(N__29461),
            .I(N__29444));
    LocalMux I__6514 (
            .O(N__29458),
            .I(N__29444));
    InMux I__6513 (
            .O(N__29457),
            .I(N__29441));
    Span4Mux_h I__6512 (
            .O(N__29452),
            .I(N__29438));
    Span4Mux_v I__6511 (
            .O(N__29449),
            .I(N__29433));
    Span4Mux_v I__6510 (
            .O(N__29444),
            .I(N__29433));
    LocalMux I__6509 (
            .O(N__29441),
            .I(N__29430));
    Span4Mux_v I__6508 (
            .O(N__29438),
            .I(N__29427));
    Span4Mux_h I__6507 (
            .O(N__29433),
            .I(N__29424));
    Span4Mux_h I__6506 (
            .O(N__29430),
            .I(N__29421));
    Odrv4 I__6505 (
            .O(N__29427),
            .I(wrtrigval_2));
    Odrv4 I__6504 (
            .O(N__29424),
            .I(wrtrigval_2));
    Odrv4 I__6503 (
            .O(N__29421),
            .I(wrtrigval_2));
    InMux I__6502 (
            .O(N__29414),
            .I(N__29410));
    InMux I__6501 (
            .O(N__29413),
            .I(N__29407));
    LocalMux I__6500 (
            .O(N__29410),
            .I(N__29404));
    LocalMux I__6499 (
            .O(N__29407),
            .I(configRegister_17));
    Odrv4 I__6498 (
            .O(N__29404),
            .I(configRegister_17));
    CascadeMux I__6497 (
            .O(N__29399),
            .I(N__29396));
    InMux I__6496 (
            .O(N__29396),
            .I(N__29391));
    InMux I__6495 (
            .O(N__29395),
            .I(N__29388));
    InMux I__6494 (
            .O(N__29394),
            .I(N__29385));
    LocalMux I__6493 (
            .O(N__29391),
            .I(N__29379));
    LocalMux I__6492 (
            .O(N__29388),
            .I(N__29374));
    LocalMux I__6491 (
            .O(N__29385),
            .I(N__29374));
    InMux I__6490 (
            .O(N__29384),
            .I(N__29369));
    InMux I__6489 (
            .O(N__29383),
            .I(N__29369));
    InMux I__6488 (
            .O(N__29382),
            .I(N__29366));
    Span4Mux_h I__6487 (
            .O(N__29379),
            .I(N__29363));
    Span4Mux_h I__6486 (
            .O(N__29374),
            .I(N__29356));
    LocalMux I__6485 (
            .O(N__29369),
            .I(N__29356));
    LocalMux I__6484 (
            .O(N__29366),
            .I(N__29356));
    Span4Mux_v I__6483 (
            .O(N__29363),
            .I(N__29351));
    Span4Mux_v I__6482 (
            .O(N__29356),
            .I(N__29348));
    InMux I__6481 (
            .O(N__29355),
            .I(N__29345));
    InMux I__6480 (
            .O(N__29354),
            .I(N__29342));
    Odrv4 I__6479 (
            .O(N__29351),
            .I(cmd_21));
    Odrv4 I__6478 (
            .O(N__29348),
            .I(cmd_21));
    LocalMux I__6477 (
            .O(N__29345),
            .I(cmd_21));
    LocalMux I__6476 (
            .O(N__29342),
            .I(cmd_21));
    InMux I__6475 (
            .O(N__29333),
            .I(N__29327));
    InMux I__6474 (
            .O(N__29332),
            .I(N__29321));
    InMux I__6473 (
            .O(N__29331),
            .I(N__29315));
    InMux I__6472 (
            .O(N__29330),
            .I(N__29312));
    LocalMux I__6471 (
            .O(N__29327),
            .I(N__29307));
    InMux I__6470 (
            .O(N__29326),
            .I(N__29304));
    InMux I__6469 (
            .O(N__29325),
            .I(N__29301));
    CascadeMux I__6468 (
            .O(N__29324),
            .I(N__29296));
    LocalMux I__6467 (
            .O(N__29321),
            .I(N__29287));
    InMux I__6466 (
            .O(N__29320),
            .I(N__29284));
    InMux I__6465 (
            .O(N__29319),
            .I(N__29279));
    InMux I__6464 (
            .O(N__29318),
            .I(N__29279));
    LocalMux I__6463 (
            .O(N__29315),
            .I(N__29274));
    LocalMux I__6462 (
            .O(N__29312),
            .I(N__29274));
    InMux I__6461 (
            .O(N__29311),
            .I(N__29271));
    InMux I__6460 (
            .O(N__29310),
            .I(N__29268));
    Span4Mux_v I__6459 (
            .O(N__29307),
            .I(N__29262));
    LocalMux I__6458 (
            .O(N__29304),
            .I(N__29262));
    LocalMux I__6457 (
            .O(N__29301),
            .I(N__29259));
    InMux I__6456 (
            .O(N__29300),
            .I(N__29254));
    InMux I__6455 (
            .O(N__29299),
            .I(N__29254));
    InMux I__6454 (
            .O(N__29296),
            .I(N__29243));
    InMux I__6453 (
            .O(N__29295),
            .I(N__29243));
    InMux I__6452 (
            .O(N__29294),
            .I(N__29243));
    InMux I__6451 (
            .O(N__29293),
            .I(N__29240));
    InMux I__6450 (
            .O(N__29292),
            .I(N__29237));
    InMux I__6449 (
            .O(N__29291),
            .I(N__29234));
    InMux I__6448 (
            .O(N__29290),
            .I(N__29231));
    Span4Mux_h I__6447 (
            .O(N__29287),
            .I(N__29224));
    LocalMux I__6446 (
            .O(N__29284),
            .I(N__29224));
    LocalMux I__6445 (
            .O(N__29279),
            .I(N__29224));
    Span4Mux_h I__6444 (
            .O(N__29274),
            .I(N__29217));
    LocalMux I__6443 (
            .O(N__29271),
            .I(N__29217));
    LocalMux I__6442 (
            .O(N__29268),
            .I(N__29217));
    InMux I__6441 (
            .O(N__29267),
            .I(N__29214));
    Span4Mux_v I__6440 (
            .O(N__29262),
            .I(N__29211));
    Span4Mux_h I__6439 (
            .O(N__29259),
            .I(N__29206));
    LocalMux I__6438 (
            .O(N__29254),
            .I(N__29206));
    InMux I__6437 (
            .O(N__29253),
            .I(N__29197));
    InMux I__6436 (
            .O(N__29252),
            .I(N__29197));
    InMux I__6435 (
            .O(N__29251),
            .I(N__29197));
    InMux I__6434 (
            .O(N__29250),
            .I(N__29197));
    LocalMux I__6433 (
            .O(N__29243),
            .I(N__29194));
    LocalMux I__6432 (
            .O(N__29240),
            .I(N__29187));
    LocalMux I__6431 (
            .O(N__29237),
            .I(N__29187));
    LocalMux I__6430 (
            .O(N__29234),
            .I(N__29187));
    LocalMux I__6429 (
            .O(N__29231),
            .I(N__29184));
    Span4Mux_v I__6428 (
            .O(N__29224),
            .I(N__29179));
    Span4Mux_v I__6427 (
            .O(N__29217),
            .I(N__29179));
    LocalMux I__6426 (
            .O(N__29214),
            .I(N__29176));
    Span4Mux_h I__6425 (
            .O(N__29211),
            .I(N__29171));
    Span4Mux_h I__6424 (
            .O(N__29206),
            .I(N__29171));
    LocalMux I__6423 (
            .O(N__29197),
            .I(N__29164));
    Span4Mux_s3_v I__6422 (
            .O(N__29194),
            .I(N__29164));
    Span4Mux_v I__6421 (
            .O(N__29187),
            .I(N__29164));
    Span4Mux_v I__6420 (
            .O(N__29184),
            .I(N__29159));
    Span4Mux_h I__6419 (
            .O(N__29179),
            .I(N__29159));
    Span4Mux_h I__6418 (
            .O(N__29176),
            .I(N__29152));
    Span4Mux_v I__6417 (
            .O(N__29171),
            .I(N__29152));
    Span4Mux_h I__6416 (
            .O(N__29164),
            .I(N__29152));
    Odrv4 I__6415 (
            .O(N__29159),
            .I(wrtrigcfg_1));
    Odrv4 I__6414 (
            .O(N__29152),
            .I(wrtrigcfg_1));
    InMux I__6413 (
            .O(N__29147),
            .I(N__29144));
    LocalMux I__6412 (
            .O(N__29144),
            .I(N__29140));
    InMux I__6411 (
            .O(N__29143),
            .I(N__29137));
    Odrv12 I__6410 (
            .O(N__29140),
            .I(configRegister_14_adj_1306));
    LocalMux I__6409 (
            .O(N__29137),
            .I(configRegister_14_adj_1306));
    InMux I__6408 (
            .O(N__29132),
            .I(N__29124));
    InMux I__6407 (
            .O(N__29131),
            .I(N__29119));
    InMux I__6406 (
            .O(N__29130),
            .I(N__29116));
    InMux I__6405 (
            .O(N__29129),
            .I(N__29111));
    CascadeMux I__6404 (
            .O(N__29128),
            .I(N__29104));
    InMux I__6403 (
            .O(N__29127),
            .I(N__29101));
    LocalMux I__6402 (
            .O(N__29124),
            .I(N__29098));
    InMux I__6401 (
            .O(N__29123),
            .I(N__29092));
    InMux I__6400 (
            .O(N__29122),
            .I(N__29092));
    LocalMux I__6399 (
            .O(N__29119),
            .I(N__29089));
    LocalMux I__6398 (
            .O(N__29116),
            .I(N__29086));
    InMux I__6397 (
            .O(N__29115),
            .I(N__29083));
    InMux I__6396 (
            .O(N__29114),
            .I(N__29080));
    LocalMux I__6395 (
            .O(N__29111),
            .I(N__29077));
    InMux I__6394 (
            .O(N__29110),
            .I(N__29074));
    InMux I__6393 (
            .O(N__29109),
            .I(N__29071));
    InMux I__6392 (
            .O(N__29108),
            .I(N__29068));
    InMux I__6391 (
            .O(N__29107),
            .I(N__29065));
    InMux I__6390 (
            .O(N__29104),
            .I(N__29060));
    LocalMux I__6389 (
            .O(N__29101),
            .I(N__29057));
    Span4Mux_h I__6388 (
            .O(N__29098),
            .I(N__29054));
    InMux I__6387 (
            .O(N__29097),
            .I(N__29051));
    LocalMux I__6386 (
            .O(N__29092),
            .I(N__29044));
    Span4Mux_v I__6385 (
            .O(N__29089),
            .I(N__29044));
    Span4Mux_v I__6384 (
            .O(N__29086),
            .I(N__29044));
    LocalMux I__6383 (
            .O(N__29083),
            .I(N__29041));
    LocalMux I__6382 (
            .O(N__29080),
            .I(N__29036));
    Span4Mux_v I__6381 (
            .O(N__29077),
            .I(N__29036));
    LocalMux I__6380 (
            .O(N__29074),
            .I(N__29027));
    LocalMux I__6379 (
            .O(N__29071),
            .I(N__29027));
    LocalMux I__6378 (
            .O(N__29068),
            .I(N__29027));
    LocalMux I__6377 (
            .O(N__29065),
            .I(N__29027));
    InMux I__6376 (
            .O(N__29064),
            .I(N__29024));
    InMux I__6375 (
            .O(N__29063),
            .I(N__29021));
    LocalMux I__6374 (
            .O(N__29060),
            .I(N__29018));
    Span4Mux_h I__6373 (
            .O(N__29057),
            .I(N__29015));
    Span4Mux_v I__6372 (
            .O(N__29054),
            .I(N__29012));
    LocalMux I__6371 (
            .O(N__29051),
            .I(N__29007));
    Span4Mux_h I__6370 (
            .O(N__29044),
            .I(N__29007));
    Span4Mux_v I__6369 (
            .O(N__29041),
            .I(N__29000));
    Span4Mux_h I__6368 (
            .O(N__29036),
            .I(N__29000));
    Span4Mux_v I__6367 (
            .O(N__29027),
            .I(N__29000));
    LocalMux I__6366 (
            .O(N__29024),
            .I(cmd_12));
    LocalMux I__6365 (
            .O(N__29021),
            .I(cmd_12));
    Odrv12 I__6364 (
            .O(N__29018),
            .I(cmd_12));
    Odrv4 I__6363 (
            .O(N__29015),
            .I(cmd_12));
    Odrv4 I__6362 (
            .O(N__29012),
            .I(cmd_12));
    Odrv4 I__6361 (
            .O(N__29007),
            .I(cmd_12));
    Odrv4 I__6360 (
            .O(N__29000),
            .I(cmd_12));
    CascadeMux I__6359 (
            .O(N__28985),
            .I(N__28982));
    InMux I__6358 (
            .O(N__28982),
            .I(N__28979));
    LocalMux I__6357 (
            .O(N__28979),
            .I(N__28975));
    InMux I__6356 (
            .O(N__28978),
            .I(N__28972));
    Span4Mux_h I__6355 (
            .O(N__28975),
            .I(N__28969));
    LocalMux I__6354 (
            .O(N__28972),
            .I(fwd_7));
    Odrv4 I__6353 (
            .O(N__28969),
            .I(fwd_7));
    InMux I__6352 (
            .O(N__28964),
            .I(N__28958));
    InMux I__6351 (
            .O(N__28963),
            .I(N__28958));
    LocalMux I__6350 (
            .O(N__28958),
            .I(N__28951));
    InMux I__6349 (
            .O(N__28957),
            .I(N__28946));
    InMux I__6348 (
            .O(N__28956),
            .I(N__28946));
    InMux I__6347 (
            .O(N__28955),
            .I(N__28941));
    InMux I__6346 (
            .O(N__28954),
            .I(N__28941));
    Span4Mux_v I__6345 (
            .O(N__28951),
            .I(N__28938));
    LocalMux I__6344 (
            .O(N__28946),
            .I(N__28935));
    LocalMux I__6343 (
            .O(N__28941),
            .I(\Inst_core.Inst_trigger.levelReg_0 ));
    Odrv4 I__6342 (
            .O(N__28938),
            .I(\Inst_core.Inst_trigger.levelReg_0 ));
    Odrv4 I__6341 (
            .O(N__28935),
            .I(\Inst_core.Inst_trigger.levelReg_0 ));
    InMux I__6340 (
            .O(N__28928),
            .I(N__28924));
    InMux I__6339 (
            .O(N__28927),
            .I(N__28921));
    LocalMux I__6338 (
            .O(N__28924),
            .I(N__28918));
    LocalMux I__6337 (
            .O(N__28921),
            .I(configRegister_17_adj_1343));
    Odrv4 I__6336 (
            .O(N__28918),
            .I(configRegister_17_adj_1343));
    InMux I__6335 (
            .O(N__28913),
            .I(N__28904));
    InMux I__6334 (
            .O(N__28912),
            .I(N__28904));
    InMux I__6333 (
            .O(N__28911),
            .I(N__28899));
    InMux I__6332 (
            .O(N__28910),
            .I(N__28899));
    InMux I__6331 (
            .O(N__28909),
            .I(N__28896));
    LocalMux I__6330 (
            .O(N__28904),
            .I(N__28893));
    LocalMux I__6329 (
            .O(N__28899),
            .I(N__28890));
    LocalMux I__6328 (
            .O(N__28896),
            .I(N__28885));
    Span4Mux_v I__6327 (
            .O(N__28893),
            .I(N__28885));
    Odrv4 I__6326 (
            .O(N__28890),
            .I(\Inst_core.Inst_trigger.levelReg_1 ));
    Odrv4 I__6325 (
            .O(N__28885),
            .I(\Inst_core.Inst_trigger.levelReg_1 ));
    InMux I__6324 (
            .O(N__28880),
            .I(N__28874));
    InMux I__6323 (
            .O(N__28879),
            .I(N__28874));
    LocalMux I__6322 (
            .O(N__28874),
            .I(N__28871));
    Span12Mux_s5_v I__6321 (
            .O(N__28871),
            .I(N__28868));
    Odrv12 I__6320 (
            .O(N__28868),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n99 ));
    InMux I__6319 (
            .O(N__28865),
            .I(N__28862));
    LocalMux I__6318 (
            .O(N__28862),
            .I(N__28858));
    InMux I__6317 (
            .O(N__28861),
            .I(N__28855));
    Odrv12 I__6316 (
            .O(N__28858),
            .I(valueRegister_4_adj_1372));
    LocalMux I__6315 (
            .O(N__28855),
            .I(valueRegister_4_adj_1372));
    CascadeMux I__6314 (
            .O(N__28850),
            .I(N__28847));
    InMux I__6313 (
            .O(N__28847),
            .I(N__28844));
    LocalMux I__6312 (
            .O(N__28844),
            .I(N__28840));
    InMux I__6311 (
            .O(N__28843),
            .I(N__28837));
    Odrv12 I__6310 (
            .O(N__28840),
            .I(configRegister_15_adj_1305));
    LocalMux I__6309 (
            .O(N__28837),
            .I(configRegister_15_adj_1305));
    CascadeMux I__6308 (
            .O(N__28832),
            .I(N__28829));
    InMux I__6307 (
            .O(N__28829),
            .I(N__28826));
    LocalMux I__6306 (
            .O(N__28826),
            .I(N__28822));
    InMux I__6305 (
            .O(N__28825),
            .I(N__28819));
    Span4Mux_h I__6304 (
            .O(N__28822),
            .I(N__28816));
    LocalMux I__6303 (
            .O(N__28819),
            .I(bwd_15));
    Odrv4 I__6302 (
            .O(N__28816),
            .I(bwd_15));
    InMux I__6301 (
            .O(N__28811),
            .I(N__28808));
    LocalMux I__6300 (
            .O(N__28808),
            .I(N__28805));
    Span4Mux_v I__6299 (
            .O(N__28805),
            .I(N__28801));
    InMux I__6298 (
            .O(N__28804),
            .I(N__28798));
    Odrv4 I__6297 (
            .O(N__28801),
            .I(configRegister_13_adj_1307));
    LocalMux I__6296 (
            .O(N__28798),
            .I(configRegister_13_adj_1307));
    InMux I__6295 (
            .O(N__28793),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7896 ));
    CascadeMux I__6294 (
            .O(N__28790),
            .I(N__28786));
    InMux I__6293 (
            .O(N__28789),
            .I(N__28783));
    InMux I__6292 (
            .O(N__28786),
            .I(N__28780));
    LocalMux I__6291 (
            .O(N__28783),
            .I(N__28777));
    LocalMux I__6290 (
            .O(N__28780),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14 ));
    Odrv4 I__6289 (
            .O(N__28777),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14 ));
    InMux I__6288 (
            .O(N__28772),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7897 ));
    InMux I__6287 (
            .O(N__28769),
            .I(N__28763));
    CascadeMux I__6286 (
            .O(N__28768),
            .I(N__28758));
    CascadeMux I__6285 (
            .O(N__28767),
            .I(N__28754));
    CascadeMux I__6284 (
            .O(N__28766),
            .I(N__28750));
    LocalMux I__6283 (
            .O(N__28763),
            .I(N__28746));
    InMux I__6282 (
            .O(N__28762),
            .I(N__28726));
    InMux I__6281 (
            .O(N__28761),
            .I(N__28726));
    InMux I__6280 (
            .O(N__28758),
            .I(N__28726));
    InMux I__6279 (
            .O(N__28757),
            .I(N__28726));
    InMux I__6278 (
            .O(N__28754),
            .I(N__28726));
    InMux I__6277 (
            .O(N__28753),
            .I(N__28726));
    InMux I__6276 (
            .O(N__28750),
            .I(N__28726));
    InMux I__6275 (
            .O(N__28749),
            .I(N__28726));
    Span4Mux_h I__6274 (
            .O(N__28746),
            .I(N__28723));
    CascadeMux I__6273 (
            .O(N__28745),
            .I(N__28719));
    CascadeMux I__6272 (
            .O(N__28744),
            .I(N__28715));
    CascadeMux I__6271 (
            .O(N__28743),
            .I(N__28711));
    LocalMux I__6270 (
            .O(N__28726),
            .I(N__28705));
    Span4Mux_v I__6269 (
            .O(N__28723),
            .I(N__28705));
    InMux I__6268 (
            .O(N__28722),
            .I(N__28690));
    InMux I__6267 (
            .O(N__28719),
            .I(N__28690));
    InMux I__6266 (
            .O(N__28718),
            .I(N__28690));
    InMux I__6265 (
            .O(N__28715),
            .I(N__28690));
    InMux I__6264 (
            .O(N__28714),
            .I(N__28690));
    InMux I__6263 (
            .O(N__28711),
            .I(N__28690));
    InMux I__6262 (
            .O(N__28710),
            .I(N__28690));
    Span4Mux_v I__6261 (
            .O(N__28705),
            .I(N__28687));
    LocalMux I__6260 (
            .O(N__28690),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n1662 ));
    Odrv4 I__6259 (
            .O(N__28687),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n1662 ));
    InMux I__6258 (
            .O(N__28682),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7898 ));
    CascadeMux I__6257 (
            .O(N__28679),
            .I(N__28676));
    InMux I__6256 (
            .O(N__28676),
            .I(N__28672));
    InMux I__6255 (
            .O(N__28675),
            .I(N__28669));
    LocalMux I__6254 (
            .O(N__28672),
            .I(N__28666));
    LocalMux I__6253 (
            .O(N__28669),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15 ));
    Odrv4 I__6252 (
            .O(N__28666),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15 ));
    CEMux I__6251 (
            .O(N__28661),
            .I(N__28658));
    LocalMux I__6250 (
            .O(N__28658),
            .I(N__28654));
    CEMux I__6249 (
            .O(N__28657),
            .I(N__28651));
    Odrv12 I__6248 (
            .O(N__28654),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4144 ));
    LocalMux I__6247 (
            .O(N__28651),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4144 ));
    InMux I__6246 (
            .O(N__28646),
            .I(N__28643));
    LocalMux I__6245 (
            .O(N__28643),
            .I(N__28639));
    CascadeMux I__6244 (
            .O(N__28642),
            .I(N__28636));
    Span4Mux_v I__6243 (
            .O(N__28639),
            .I(N__28632));
    InMux I__6242 (
            .O(N__28636),
            .I(N__28627));
    InMux I__6241 (
            .O(N__28635),
            .I(N__28627));
    Odrv4 I__6240 (
            .O(N__28632),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2 ));
    LocalMux I__6239 (
            .O(N__28627),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2 ));
    SRMux I__6238 (
            .O(N__28622),
            .I(N__28619));
    LocalMux I__6237 (
            .O(N__28619),
            .I(N__28616));
    Span4Mux_s2_h I__6236 (
            .O(N__28616),
            .I(N__28613));
    Span4Mux_h I__6235 (
            .O(N__28613),
            .I(N__28610));
    Odrv4 I__6234 (
            .O(N__28610),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4761 ));
    CascadeMux I__6233 (
            .O(N__28607),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n2_cascade_ ));
    InMux I__6232 (
            .O(N__28604),
            .I(N__28601));
    LocalMux I__6231 (
            .O(N__28601),
            .I(N__28598));
    Span4Mux_v I__6230 (
            .O(N__28598),
            .I(N__28595));
    Sp12to4 I__6229 (
            .O(N__28595),
            .I(N__28592));
    Odrv12 I__6228 (
            .O(N__28592),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register ));
    InMux I__6227 (
            .O(N__28589),
            .I(N__28586));
    LocalMux I__6226 (
            .O(N__28586),
            .I(N__28583));
    Span4Mux_v I__6225 (
            .O(N__28583),
            .I(N__28580));
    Odrv4 I__6224 (
            .O(N__28580),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n100 ));
    CascadeMux I__6223 (
            .O(N__28577),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n100_cascade_ ));
    InMux I__6222 (
            .O(N__28574),
            .I(N__28570));
    CascadeMux I__6221 (
            .O(N__28573),
            .I(N__28567));
    LocalMux I__6220 (
            .O(N__28570),
            .I(N__28564));
    InMux I__6219 (
            .O(N__28567),
            .I(N__28561));
    Span4Mux_s2_h I__6218 (
            .O(N__28564),
            .I(N__28558));
    LocalMux I__6217 (
            .O(N__28561),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n450 ));
    Odrv4 I__6216 (
            .O(N__28558),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n450 ));
    InMux I__6215 (
            .O(N__28553),
            .I(N__28550));
    LocalMux I__6214 (
            .O(N__28550),
            .I(N__28546));
    InMux I__6213 (
            .O(N__28549),
            .I(N__28543));
    Odrv4 I__6212 (
            .O(N__28546),
            .I(configRegister_5_adj_1315));
    LocalMux I__6211 (
            .O(N__28543),
            .I(configRegister_5_adj_1315));
    InMux I__6210 (
            .O(N__28538),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7888 ));
    InMux I__6209 (
            .O(N__28535),
            .I(N__28532));
    LocalMux I__6208 (
            .O(N__28532),
            .I(N__28528));
    InMux I__6207 (
            .O(N__28531),
            .I(N__28525));
    Odrv4 I__6206 (
            .O(N__28528),
            .I(configRegister_6_adj_1314));
    LocalMux I__6205 (
            .O(N__28525),
            .I(configRegister_6_adj_1314));
    InMux I__6204 (
            .O(N__28520),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7889 ));
    InMux I__6203 (
            .O(N__28517),
            .I(N__28514));
    LocalMux I__6202 (
            .O(N__28514),
            .I(N__28511));
    Span4Mux_v I__6201 (
            .O(N__28511),
            .I(N__28508));
    Span4Mux_s1_h I__6200 (
            .O(N__28508),
            .I(N__28504));
    InMux I__6199 (
            .O(N__28507),
            .I(N__28501));
    Odrv4 I__6198 (
            .O(N__28504),
            .I(configRegister_7_adj_1313));
    LocalMux I__6197 (
            .O(N__28501),
            .I(configRegister_7_adj_1313));
    InMux I__6196 (
            .O(N__28496),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7890 ));
    InMux I__6195 (
            .O(N__28493),
            .I(N__28490));
    LocalMux I__6194 (
            .O(N__28490),
            .I(N__28486));
    CascadeMux I__6193 (
            .O(N__28489),
            .I(N__28483));
    Span12Mux_s5_h I__6192 (
            .O(N__28486),
            .I(N__28480));
    InMux I__6191 (
            .O(N__28483),
            .I(N__28477));
    Odrv12 I__6190 (
            .O(N__28480),
            .I(configRegister_8_adj_1312));
    LocalMux I__6189 (
            .O(N__28477),
            .I(configRegister_8_adj_1312));
    InMux I__6188 (
            .O(N__28472),
            .I(bfn_11_5_0_));
    InMux I__6187 (
            .O(N__28469),
            .I(N__28466));
    LocalMux I__6186 (
            .O(N__28466),
            .I(N__28463));
    Span4Mux_s2_h I__6185 (
            .O(N__28463),
            .I(N__28459));
    InMux I__6184 (
            .O(N__28462),
            .I(N__28456));
    Odrv4 I__6183 (
            .O(N__28459),
            .I(configRegister_9_adj_1311));
    LocalMux I__6182 (
            .O(N__28456),
            .I(configRegister_9_adj_1311));
    InMux I__6181 (
            .O(N__28451),
            .I(N__28447));
    InMux I__6180 (
            .O(N__28450),
            .I(N__28444));
    LocalMux I__6179 (
            .O(N__28447),
            .I(N__28441));
    LocalMux I__6178 (
            .O(N__28444),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9 ));
    Odrv4 I__6177 (
            .O(N__28441),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9 ));
    InMux I__6176 (
            .O(N__28436),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7892 ));
    InMux I__6175 (
            .O(N__28433),
            .I(N__28430));
    LocalMux I__6174 (
            .O(N__28430),
            .I(N__28427));
    Span4Mux_v I__6173 (
            .O(N__28427),
            .I(N__28423));
    InMux I__6172 (
            .O(N__28426),
            .I(N__28420));
    Odrv4 I__6171 (
            .O(N__28423),
            .I(configRegister_10_adj_1310));
    LocalMux I__6170 (
            .O(N__28420),
            .I(configRegister_10_adj_1310));
    InMux I__6169 (
            .O(N__28415),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7893 ));
    InMux I__6168 (
            .O(N__28412),
            .I(N__28409));
    LocalMux I__6167 (
            .O(N__28409),
            .I(N__28406));
    Span4Mux_h I__6166 (
            .O(N__28406),
            .I(N__28402));
    InMux I__6165 (
            .O(N__28405),
            .I(N__28399));
    Odrv4 I__6164 (
            .O(N__28402),
            .I(configRegister_11_adj_1309));
    LocalMux I__6163 (
            .O(N__28399),
            .I(configRegister_11_adj_1309));
    InMux I__6162 (
            .O(N__28394),
            .I(N__28390));
    InMux I__6161 (
            .O(N__28393),
            .I(N__28387));
    LocalMux I__6160 (
            .O(N__28390),
            .I(N__28384));
    LocalMux I__6159 (
            .O(N__28387),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11 ));
    Odrv4 I__6158 (
            .O(N__28384),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11 ));
    InMux I__6157 (
            .O(N__28379),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7894 ));
    InMux I__6156 (
            .O(N__28376),
            .I(N__28373));
    LocalMux I__6155 (
            .O(N__28373),
            .I(N__28369));
    InMux I__6154 (
            .O(N__28372),
            .I(N__28366));
    Odrv12 I__6153 (
            .O(N__28369),
            .I(configRegister_12_adj_1308));
    LocalMux I__6152 (
            .O(N__28366),
            .I(configRegister_12_adj_1308));
    InMux I__6151 (
            .O(N__28361),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7895 ));
    InMux I__6150 (
            .O(N__28358),
            .I(N__28355));
    LocalMux I__6149 (
            .O(N__28355),
            .I(N__28352));
    Span4Mux_s2_v I__6148 (
            .O(N__28352),
            .I(N__28348));
    InMux I__6147 (
            .O(N__28351),
            .I(N__28345));
    Odrv4 I__6146 (
            .O(N__28348),
            .I(\Inst_core.n8837 ));
    LocalMux I__6145 (
            .O(N__28345),
            .I(\Inst_core.n8837 ));
    InMux I__6144 (
            .O(N__28340),
            .I(N__28334));
    InMux I__6143 (
            .O(N__28339),
            .I(N__28327));
    InMux I__6142 (
            .O(N__28338),
            .I(N__28327));
    InMux I__6141 (
            .O(N__28337),
            .I(N__28327));
    LocalMux I__6140 (
            .O(N__28334),
            .I(N__28321));
    LocalMux I__6139 (
            .O(N__28327),
            .I(N__28321));
    InMux I__6138 (
            .O(N__28326),
            .I(N__28318));
    Span4Mux_v I__6137 (
            .O(N__28321),
            .I(N__28315));
    LocalMux I__6136 (
            .O(N__28318),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.state_1 ));
    Odrv4 I__6135 (
            .O(N__28315),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.state_1 ));
    InMux I__6134 (
            .O(N__28310),
            .I(N__28306));
    InMux I__6133 (
            .O(N__28309),
            .I(N__28303));
    LocalMux I__6132 (
            .O(N__28306),
            .I(N__28300));
    LocalMux I__6131 (
            .O(N__28303),
            .I(configRegister_0_adj_1320));
    Odrv4 I__6130 (
            .O(N__28300),
            .I(configRegister_0_adj_1320));
    InMux I__6129 (
            .O(N__28295),
            .I(N__28292));
    LocalMux I__6128 (
            .O(N__28292),
            .I(N__28289));
    Span4Mux_s2_h I__6127 (
            .O(N__28289),
            .I(N__28286));
    Span4Mux_v I__6126 (
            .O(N__28286),
            .I(N__28283));
    Odrv4 I__6125 (
            .O(N__28283),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9055 ));
    InMux I__6124 (
            .O(N__28280),
            .I(bfn_11_4_0_));
    InMux I__6123 (
            .O(N__28277),
            .I(N__28274));
    LocalMux I__6122 (
            .O(N__28274),
            .I(N__28271));
    Span4Mux_s1_h I__6121 (
            .O(N__28271),
            .I(N__28267));
    InMux I__6120 (
            .O(N__28270),
            .I(N__28264));
    Odrv4 I__6119 (
            .O(N__28267),
            .I(configRegister_1_adj_1319));
    LocalMux I__6118 (
            .O(N__28264),
            .I(configRegister_1_adj_1319));
    InMux I__6117 (
            .O(N__28259),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7884 ));
    InMux I__6116 (
            .O(N__28256),
            .I(N__28252));
    InMux I__6115 (
            .O(N__28255),
            .I(N__28249));
    LocalMux I__6114 (
            .O(N__28252),
            .I(N__28246));
    LocalMux I__6113 (
            .O(N__28249),
            .I(configRegister_2_adj_1318));
    Odrv4 I__6112 (
            .O(N__28246),
            .I(configRegister_2_adj_1318));
    InMux I__6111 (
            .O(N__28241),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7885 ));
    InMux I__6110 (
            .O(N__28238),
            .I(N__28235));
    LocalMux I__6109 (
            .O(N__28235),
            .I(N__28231));
    InMux I__6108 (
            .O(N__28234),
            .I(N__28228));
    Odrv4 I__6107 (
            .O(N__28231),
            .I(configRegister_3_adj_1317));
    LocalMux I__6106 (
            .O(N__28228),
            .I(configRegister_3_adj_1317));
    InMux I__6105 (
            .O(N__28223),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7886 ));
    InMux I__6104 (
            .O(N__28220),
            .I(N__28217));
    LocalMux I__6103 (
            .O(N__28217),
            .I(N__28214));
    Span4Mux_s3_h I__6102 (
            .O(N__28214),
            .I(N__28210));
    InMux I__6101 (
            .O(N__28213),
            .I(N__28207));
    Odrv4 I__6100 (
            .O(N__28210),
            .I(configRegister_4_adj_1316));
    LocalMux I__6099 (
            .O(N__28207),
            .I(configRegister_4_adj_1316));
    InMux I__6098 (
            .O(N__28202),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7887 ));
    InMux I__6097 (
            .O(N__28199),
            .I(N__28196));
    LocalMux I__6096 (
            .O(N__28196),
            .I(N__28193));
    Span4Mux_s3_v I__6095 (
            .O(N__28193),
            .I(N__28187));
    InMux I__6094 (
            .O(N__28192),
            .I(N__28184));
    InMux I__6093 (
            .O(N__28191),
            .I(N__28179));
    InMux I__6092 (
            .O(N__28190),
            .I(N__28179));
    Span4Mux_h I__6091 (
            .O(N__28187),
            .I(N__28171));
    LocalMux I__6090 (
            .O(N__28184),
            .I(N__28171));
    LocalMux I__6089 (
            .O(N__28179),
            .I(N__28168));
    InMux I__6088 (
            .O(N__28178),
            .I(N__28165));
    InMux I__6087 (
            .O(N__28177),
            .I(N__28162));
    CascadeMux I__6086 (
            .O(N__28176),
            .I(N__28159));
    Span4Mux_v I__6085 (
            .O(N__28171),
            .I(N__28156));
    Span12Mux_s4_h I__6084 (
            .O(N__28168),
            .I(N__28151));
    LocalMux I__6083 (
            .O(N__28165),
            .I(N__28151));
    LocalMux I__6082 (
            .O(N__28162),
            .I(N__28148));
    InMux I__6081 (
            .O(N__28159),
            .I(N__28145));
    Odrv4 I__6080 (
            .O(N__28156),
            .I(cmd_35));
    Odrv12 I__6079 (
            .O(N__28151),
            .I(cmd_35));
    Odrv4 I__6078 (
            .O(N__28148),
            .I(cmd_35));
    LocalMux I__6077 (
            .O(N__28145),
            .I(cmd_35));
    InMux I__6076 (
            .O(N__28136),
            .I(N__28133));
    LocalMux I__6075 (
            .O(N__28133),
            .I(N__28129));
    InMux I__6074 (
            .O(N__28132),
            .I(N__28126));
    Odrv4 I__6073 (
            .O(N__28129),
            .I(configRegister_0_adj_1360));
    LocalMux I__6072 (
            .O(N__28126),
            .I(configRegister_0_adj_1360));
    InMux I__6071 (
            .O(N__28121),
            .I(N__28117));
    CascadeMux I__6070 (
            .O(N__28120),
            .I(N__28114));
    LocalMux I__6069 (
            .O(N__28117),
            .I(N__28110));
    InMux I__6068 (
            .O(N__28114),
            .I(N__28105));
    InMux I__6067 (
            .O(N__28113),
            .I(N__28105));
    Span4Mux_h I__6066 (
            .O(N__28110),
            .I(N__28102));
    LocalMux I__6065 (
            .O(N__28105),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4 ));
    Odrv4 I__6064 (
            .O(N__28102),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4 ));
    CascadeMux I__6063 (
            .O(N__28097),
            .I(N__28094));
    InMux I__6062 (
            .O(N__28094),
            .I(N__28091));
    LocalMux I__6061 (
            .O(N__28091),
            .I(N__28088));
    Span4Mux_s3_h I__6060 (
            .O(N__28088),
            .I(N__28082));
    InMux I__6059 (
            .O(N__28087),
            .I(N__28078));
    CascadeMux I__6058 (
            .O(N__28086),
            .I(N__28073));
    InMux I__6057 (
            .O(N__28085),
            .I(N__28069));
    Span4Mux_h I__6056 (
            .O(N__28082),
            .I(N__28066));
    InMux I__6055 (
            .O(N__28081),
            .I(N__28063));
    LocalMux I__6054 (
            .O(N__28078),
            .I(N__28060));
    InMux I__6053 (
            .O(N__28077),
            .I(N__28057));
    InMux I__6052 (
            .O(N__28076),
            .I(N__28054));
    InMux I__6051 (
            .O(N__28073),
            .I(N__28051));
    InMux I__6050 (
            .O(N__28072),
            .I(N__28048));
    LocalMux I__6049 (
            .O(N__28069),
            .I(N__28045));
    Span4Mux_v I__6048 (
            .O(N__28066),
            .I(N__28040));
    LocalMux I__6047 (
            .O(N__28063),
            .I(N__28040));
    Span4Mux_v I__6046 (
            .O(N__28060),
            .I(N__28037));
    LocalMux I__6045 (
            .O(N__28057),
            .I(N__28034));
    LocalMux I__6044 (
            .O(N__28054),
            .I(N__28029));
    LocalMux I__6043 (
            .O(N__28051),
            .I(N__28029));
    LocalMux I__6042 (
            .O(N__28048),
            .I(N__28024));
    Span4Mux_h I__6041 (
            .O(N__28045),
            .I(N__28019));
    Span4Mux_v I__6040 (
            .O(N__28040),
            .I(N__28019));
    Span4Mux_h I__6039 (
            .O(N__28037),
            .I(N__28012));
    Span4Mux_h I__6038 (
            .O(N__28034),
            .I(N__28012));
    Span4Mux_h I__6037 (
            .O(N__28029),
            .I(N__28012));
    InMux I__6036 (
            .O(N__28028),
            .I(N__28009));
    InMux I__6035 (
            .O(N__28027),
            .I(N__28006));
    Span4Mux_v I__6034 (
            .O(N__28024),
            .I(N__28001));
    Span4Mux_v I__6033 (
            .O(N__28019),
            .I(N__28001));
    Span4Mux_v I__6032 (
            .O(N__28012),
            .I(N__27998));
    LocalMux I__6031 (
            .O(N__28009),
            .I(N__27995));
    LocalMux I__6030 (
            .O(N__28006),
            .I(memoryOut_4));
    Odrv4 I__6029 (
            .O(N__28001),
            .I(memoryOut_4));
    Odrv4 I__6028 (
            .O(N__27998),
            .I(memoryOut_4));
    Odrv12 I__6027 (
            .O(N__27995),
            .I(memoryOut_4));
    SRMux I__6026 (
            .O(N__27986),
            .I(N__27983));
    LocalMux I__6025 (
            .O(N__27983),
            .I(N__27980));
    Span4Mux_s3_v I__6024 (
            .O(N__27980),
            .I(N__27977));
    Span4Mux_s1_h I__6023 (
            .O(N__27977),
            .I(N__27974));
    Span4Mux_h I__6022 (
            .O(N__27974),
            .I(N__27971));
    Odrv4 I__6021 (
            .O(N__27971),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4763 ));
    InMux I__6020 (
            .O(N__27968),
            .I(N__27965));
    LocalMux I__6019 (
            .O(N__27965),
            .I(N__27962));
    Span4Mux_s2_h I__6018 (
            .O(N__27962),
            .I(N__27959));
    Odrv4 I__6017 (
            .O(N__27959),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_5 ));
    InMux I__6016 (
            .O(N__27956),
            .I(N__27953));
    LocalMux I__6015 (
            .O(N__27953),
            .I(N__27950));
    Odrv12 I__6014 (
            .O(N__27950),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_7 ));
    CascadeMux I__6013 (
            .O(N__27947),
            .I(N__27944));
    InMux I__6012 (
            .O(N__27944),
            .I(N__27941));
    LocalMux I__6011 (
            .O(N__27941),
            .I(N__27938));
    Span4Mux_h I__6010 (
            .O(N__27938),
            .I(N__27935));
    Odrv4 I__6009 (
            .O(N__27935),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_6 ));
    InMux I__6008 (
            .O(N__27932),
            .I(N__27929));
    LocalMux I__6007 (
            .O(N__27929),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_4 ));
    InMux I__6006 (
            .O(N__27926),
            .I(N__27923));
    LocalMux I__6005 (
            .O(N__27923),
            .I(N__27920));
    Span4Mux_h I__6004 (
            .O(N__27920),
            .I(N__27917));
    Odrv4 I__6003 (
            .O(N__27917),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n11 ));
    CascadeMux I__6002 (
            .O(N__27914),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n6675_cascade_ ));
    CascadeMux I__6001 (
            .O(N__27911),
            .I(N__27907));
    InMux I__6000 (
            .O(N__27910),
            .I(N__27904));
    InMux I__5999 (
            .O(N__27907),
            .I(N__27901));
    LocalMux I__5998 (
            .O(N__27904),
            .I(N__27898));
    LocalMux I__5997 (
            .O(N__27901),
            .I(N__27895));
    Span4Mux_v I__5996 (
            .O(N__27898),
            .I(N__27892));
    Odrv4 I__5995 (
            .O(N__27895),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n564 ));
    Odrv4 I__5994 (
            .O(N__27892),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n564 ));
    CascadeMux I__5993 (
            .O(N__27887),
            .I(N__27884));
    InMux I__5992 (
            .O(N__27884),
            .I(N__27881));
    LocalMux I__5991 (
            .O(N__27881),
            .I(N__27877));
    InMux I__5990 (
            .O(N__27880),
            .I(N__27873));
    Span4Mux_v I__5989 (
            .O(N__27877),
            .I(N__27870));
    InMux I__5988 (
            .O(N__27876),
            .I(N__27867));
    LocalMux I__5987 (
            .O(N__27873),
            .I(\Inst_core.Inst_sampler.counter_17 ));
    Odrv4 I__5986 (
            .O(N__27870),
            .I(\Inst_core.Inst_sampler.counter_17 ));
    LocalMux I__5985 (
            .O(N__27867),
            .I(\Inst_core.Inst_sampler.counter_17 ));
    InMux I__5984 (
            .O(N__27860),
            .I(\Inst_core.Inst_sampler.n7964 ));
    InMux I__5983 (
            .O(N__27857),
            .I(\Inst_core.Inst_sampler.n7965 ));
    InMux I__5982 (
            .O(N__27854),
            .I(N__27851));
    LocalMux I__5981 (
            .O(N__27851),
            .I(N__27846));
    InMux I__5980 (
            .O(N__27850),
            .I(N__27843));
    InMux I__5979 (
            .O(N__27849),
            .I(N__27840));
    Span4Mux_h I__5978 (
            .O(N__27846),
            .I(N__27837));
    LocalMux I__5977 (
            .O(N__27843),
            .I(N__27834));
    LocalMux I__5976 (
            .O(N__27840),
            .I(\Inst_core.Inst_sampler.counter_19 ));
    Odrv4 I__5975 (
            .O(N__27837),
            .I(\Inst_core.Inst_sampler.counter_19 ));
    Odrv4 I__5974 (
            .O(N__27834),
            .I(\Inst_core.Inst_sampler.counter_19 ));
    InMux I__5973 (
            .O(N__27827),
            .I(\Inst_core.Inst_sampler.n7966 ));
    InMux I__5972 (
            .O(N__27824),
            .I(N__27819));
    InMux I__5971 (
            .O(N__27823),
            .I(N__27814));
    InMux I__5970 (
            .O(N__27822),
            .I(N__27814));
    LocalMux I__5969 (
            .O(N__27819),
            .I(\Inst_core.Inst_sampler.counter_20 ));
    LocalMux I__5968 (
            .O(N__27814),
            .I(\Inst_core.Inst_sampler.counter_20 ));
    InMux I__5967 (
            .O(N__27809),
            .I(\Inst_core.Inst_sampler.n7967 ));
    InMux I__5966 (
            .O(N__27806),
            .I(N__27802));
    InMux I__5965 (
            .O(N__27805),
            .I(N__27799));
    LocalMux I__5964 (
            .O(N__27802),
            .I(N__27795));
    LocalMux I__5963 (
            .O(N__27799),
            .I(N__27792));
    InMux I__5962 (
            .O(N__27798),
            .I(N__27789));
    Span4Mux_v I__5961 (
            .O(N__27795),
            .I(N__27786));
    Span4Mux_v I__5960 (
            .O(N__27792),
            .I(N__27783));
    LocalMux I__5959 (
            .O(N__27789),
            .I(\Inst_core.Inst_sampler.counter_21 ));
    Odrv4 I__5958 (
            .O(N__27786),
            .I(\Inst_core.Inst_sampler.counter_21 ));
    Odrv4 I__5957 (
            .O(N__27783),
            .I(\Inst_core.Inst_sampler.counter_21 ));
    InMux I__5956 (
            .O(N__27776),
            .I(\Inst_core.Inst_sampler.n7968 ));
    InMux I__5955 (
            .O(N__27773),
            .I(\Inst_core.Inst_sampler.n7969 ));
    InMux I__5954 (
            .O(N__27770),
            .I(\Inst_core.Inst_sampler.n7970 ));
    SRMux I__5953 (
            .O(N__27767),
            .I(N__27764));
    LocalMux I__5952 (
            .O(N__27764),
            .I(N__27760));
    SRMux I__5951 (
            .O(N__27763),
            .I(N__27757));
    Span4Mux_s1_v I__5950 (
            .O(N__27760),
            .I(N__27751));
    LocalMux I__5949 (
            .O(N__27757),
            .I(N__27751));
    SRMux I__5948 (
            .O(N__27756),
            .I(N__27748));
    Span4Mux_v I__5947 (
            .O(N__27751),
            .I(N__27745));
    LocalMux I__5946 (
            .O(N__27748),
            .I(N__27742));
    Span4Mux_s3_h I__5945 (
            .O(N__27745),
            .I(N__27737));
    Span4Mux_v I__5944 (
            .O(N__27742),
            .I(N__27737));
    Span4Mux_h I__5943 (
            .O(N__27737),
            .I(N__27734));
    Span4Mux_v I__5942 (
            .O(N__27734),
            .I(N__27731));
    Odrv4 I__5941 (
            .O(N__27731),
            .I(\Inst_core.Inst_sampler.n1700 ));
    InMux I__5940 (
            .O(N__27728),
            .I(N__27725));
    LocalMux I__5939 (
            .O(N__27725),
            .I(N__27720));
    InMux I__5938 (
            .O(N__27724),
            .I(N__27715));
    InMux I__5937 (
            .O(N__27723),
            .I(N__27715));
    Odrv4 I__5936 (
            .O(N__27720),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997 ));
    LocalMux I__5935 (
            .O(N__27715),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997 ));
    SRMux I__5934 (
            .O(N__27710),
            .I(N__27707));
    LocalMux I__5933 (
            .O(N__27707),
            .I(N__27704));
    Odrv12 I__5932 (
            .O(N__27704),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n8622 ));
    InMux I__5931 (
            .O(N__27701),
            .I(N__27696));
    InMux I__5930 (
            .O(N__27700),
            .I(N__27693));
    InMux I__5929 (
            .O(N__27699),
            .I(N__27690));
    LocalMux I__5928 (
            .O(N__27696),
            .I(N__27687));
    LocalMux I__5927 (
            .O(N__27693),
            .I(\Inst_core.Inst_sampler.counter_9 ));
    LocalMux I__5926 (
            .O(N__27690),
            .I(\Inst_core.Inst_sampler.counter_9 ));
    Odrv4 I__5925 (
            .O(N__27687),
            .I(\Inst_core.Inst_sampler.counter_9 ));
    InMux I__5924 (
            .O(N__27680),
            .I(\Inst_core.Inst_sampler.n7956 ));
    InMux I__5923 (
            .O(N__27677),
            .I(N__27670));
    InMux I__5922 (
            .O(N__27676),
            .I(N__27670));
    InMux I__5921 (
            .O(N__27675),
            .I(N__27667));
    LocalMux I__5920 (
            .O(N__27670),
            .I(N__27664));
    LocalMux I__5919 (
            .O(N__27667),
            .I(\Inst_core.Inst_sampler.counter_10 ));
    Odrv4 I__5918 (
            .O(N__27664),
            .I(\Inst_core.Inst_sampler.counter_10 ));
    InMux I__5917 (
            .O(N__27659),
            .I(\Inst_core.Inst_sampler.n7957 ));
    InMux I__5916 (
            .O(N__27656),
            .I(\Inst_core.Inst_sampler.n7958 ));
    InMux I__5915 (
            .O(N__27653),
            .I(\Inst_core.Inst_sampler.n7959 ));
    InMux I__5914 (
            .O(N__27650),
            .I(N__27645));
    InMux I__5913 (
            .O(N__27649),
            .I(N__27640));
    InMux I__5912 (
            .O(N__27648),
            .I(N__27640));
    LocalMux I__5911 (
            .O(N__27645),
            .I(\Inst_core.Inst_sampler.counter_13 ));
    LocalMux I__5910 (
            .O(N__27640),
            .I(\Inst_core.Inst_sampler.counter_13 ));
    InMux I__5909 (
            .O(N__27635),
            .I(\Inst_core.Inst_sampler.n7960 ));
    InMux I__5908 (
            .O(N__27632),
            .I(N__27627));
    InMux I__5907 (
            .O(N__27631),
            .I(N__27622));
    InMux I__5906 (
            .O(N__27630),
            .I(N__27622));
    LocalMux I__5905 (
            .O(N__27627),
            .I(\Inst_core.Inst_sampler.counter_14 ));
    LocalMux I__5904 (
            .O(N__27622),
            .I(\Inst_core.Inst_sampler.counter_14 ));
    InMux I__5903 (
            .O(N__27617),
            .I(\Inst_core.Inst_sampler.n7961 ));
    InMux I__5902 (
            .O(N__27614),
            .I(N__27609));
    InMux I__5901 (
            .O(N__27613),
            .I(N__27604));
    InMux I__5900 (
            .O(N__27612),
            .I(N__27604));
    LocalMux I__5899 (
            .O(N__27609),
            .I(\Inst_core.Inst_sampler.counter_15 ));
    LocalMux I__5898 (
            .O(N__27604),
            .I(\Inst_core.Inst_sampler.counter_15 ));
    InMux I__5897 (
            .O(N__27599),
            .I(\Inst_core.Inst_sampler.n7962 ));
    CascadeMux I__5896 (
            .O(N__27596),
            .I(N__27593));
    InMux I__5895 (
            .O(N__27593),
            .I(N__27588));
    InMux I__5894 (
            .O(N__27592),
            .I(N__27585));
    InMux I__5893 (
            .O(N__27591),
            .I(N__27582));
    LocalMux I__5892 (
            .O(N__27588),
            .I(N__27579));
    LocalMux I__5891 (
            .O(N__27585),
            .I(N__27576));
    LocalMux I__5890 (
            .O(N__27582),
            .I(\Inst_core.Inst_sampler.counter_16 ));
    Odrv12 I__5889 (
            .O(N__27579),
            .I(\Inst_core.Inst_sampler.counter_16 ));
    Odrv4 I__5888 (
            .O(N__27576),
            .I(\Inst_core.Inst_sampler.counter_16 ));
    InMux I__5887 (
            .O(N__27569),
            .I(bfn_9_16_0_));
    InMux I__5886 (
            .O(N__27566),
            .I(bfn_9_14_0_));
    InMux I__5885 (
            .O(N__27563),
            .I(\Inst_core.Inst_sampler.n7948 ));
    InMux I__5884 (
            .O(N__27560),
            .I(\Inst_core.Inst_sampler.n7949 ));
    InMux I__5883 (
            .O(N__27557),
            .I(\Inst_core.Inst_sampler.n7950 ));
    InMux I__5882 (
            .O(N__27554),
            .I(N__27549));
    InMux I__5881 (
            .O(N__27553),
            .I(N__27546));
    InMux I__5880 (
            .O(N__27552),
            .I(N__27543));
    LocalMux I__5879 (
            .O(N__27549),
            .I(\Inst_core.Inst_sampler.counter_4 ));
    LocalMux I__5878 (
            .O(N__27546),
            .I(\Inst_core.Inst_sampler.counter_4 ));
    LocalMux I__5877 (
            .O(N__27543),
            .I(\Inst_core.Inst_sampler.counter_4 ));
    InMux I__5876 (
            .O(N__27536),
            .I(\Inst_core.Inst_sampler.n7951 ));
    InMux I__5875 (
            .O(N__27533),
            .I(\Inst_core.Inst_sampler.n7952 ));
    InMux I__5874 (
            .O(N__27530),
            .I(\Inst_core.Inst_sampler.n7953 ));
    InMux I__5873 (
            .O(N__27527),
            .I(N__27522));
    InMux I__5872 (
            .O(N__27526),
            .I(N__27519));
    InMux I__5871 (
            .O(N__27525),
            .I(N__27516));
    LocalMux I__5870 (
            .O(N__27522),
            .I(\Inst_core.Inst_sampler.counter_7 ));
    LocalMux I__5869 (
            .O(N__27519),
            .I(\Inst_core.Inst_sampler.counter_7 ));
    LocalMux I__5868 (
            .O(N__27516),
            .I(\Inst_core.Inst_sampler.counter_7 ));
    InMux I__5867 (
            .O(N__27509),
            .I(\Inst_core.Inst_sampler.n7954 ));
    InMux I__5866 (
            .O(N__27506),
            .I(N__27503));
    LocalMux I__5865 (
            .O(N__27503),
            .I(N__27498));
    InMux I__5864 (
            .O(N__27502),
            .I(N__27495));
    InMux I__5863 (
            .O(N__27501),
            .I(N__27492));
    Span4Mux_h I__5862 (
            .O(N__27498),
            .I(N__27489));
    LocalMux I__5861 (
            .O(N__27495),
            .I(N__27486));
    LocalMux I__5860 (
            .O(N__27492),
            .I(\Inst_core.Inst_sampler.counter_8 ));
    Odrv4 I__5859 (
            .O(N__27489),
            .I(\Inst_core.Inst_sampler.counter_8 ));
    Odrv4 I__5858 (
            .O(N__27486),
            .I(\Inst_core.Inst_sampler.counter_8 ));
    InMux I__5857 (
            .O(N__27479),
            .I(bfn_9_15_0_));
    InMux I__5856 (
            .O(N__27476),
            .I(N__27472));
    InMux I__5855 (
            .O(N__27475),
            .I(N__27469));
    LocalMux I__5854 (
            .O(N__27472),
            .I(maskRegister_1_adj_1327));
    LocalMux I__5853 (
            .O(N__27469),
            .I(maskRegister_1_adj_1327));
    SRMux I__5852 (
            .O(N__27464),
            .I(N__27461));
    LocalMux I__5851 (
            .O(N__27461),
            .I(N__27458));
    Span4Mux_v I__5850 (
            .O(N__27458),
            .I(N__27455));
    Sp12to4 I__5849 (
            .O(N__27455),
            .I(N__27452));
    Odrv12 I__5848 (
            .O(N__27452),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4753 ));
    InMux I__5847 (
            .O(N__27449),
            .I(N__27445));
    InMux I__5846 (
            .O(N__27448),
            .I(N__27442));
    LocalMux I__5845 (
            .O(N__27445),
            .I(maskRegister_2_adj_1326));
    LocalMux I__5844 (
            .O(N__27442),
            .I(maskRegister_2_adj_1326));
    InMux I__5843 (
            .O(N__27437),
            .I(N__27433));
    InMux I__5842 (
            .O(N__27436),
            .I(N__27430));
    LocalMux I__5841 (
            .O(N__27433),
            .I(N__27427));
    LocalMux I__5840 (
            .O(N__27430),
            .I(maskRegister_3_adj_1325));
    Odrv4 I__5839 (
            .O(N__27427),
            .I(maskRegister_3_adj_1325));
    InMux I__5838 (
            .O(N__27422),
            .I(N__27419));
    LocalMux I__5837 (
            .O(N__27419),
            .I(N__27416));
    Span4Mux_s3_h I__5836 (
            .O(N__27416),
            .I(N__27412));
    InMux I__5835 (
            .O(N__27415),
            .I(N__27409));
    Odrv4 I__5834 (
            .O(N__27412),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6 ));
    LocalMux I__5833 (
            .O(N__27409),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6 ));
    InMux I__5832 (
            .O(N__27404),
            .I(N__27401));
    LocalMux I__5831 (
            .O(N__27401),
            .I(N__27398));
    Span4Mux_v I__5830 (
            .O(N__27398),
            .I(N__27395));
    Span4Mux_v I__5829 (
            .O(N__27395),
            .I(N__27391));
    InMux I__5828 (
            .O(N__27394),
            .I(N__27388));
    Odrv4 I__5827 (
            .O(N__27391),
            .I(valueRegister_6_adj_1330));
    LocalMux I__5826 (
            .O(N__27388),
            .I(valueRegister_6_adj_1330));
    InMux I__5825 (
            .O(N__27383),
            .I(N__27380));
    LocalMux I__5824 (
            .O(N__27380),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_6 ));
    SRMux I__5823 (
            .O(N__27377),
            .I(N__27374));
    LocalMux I__5822 (
            .O(N__27374),
            .I(N__27371));
    Span4Mux_v I__5821 (
            .O(N__27371),
            .I(N__27368));
    Span4Mux_s2_h I__5820 (
            .O(N__27368),
            .I(N__27365));
    Odrv4 I__5819 (
            .O(N__27365),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4758 ));
    InMux I__5818 (
            .O(N__27362),
            .I(N__27357));
    CascadeMux I__5817 (
            .O(N__27361),
            .I(N__27354));
    InMux I__5816 (
            .O(N__27360),
            .I(N__27351));
    LocalMux I__5815 (
            .O(N__27357),
            .I(N__27348));
    InMux I__5814 (
            .O(N__27354),
            .I(N__27345));
    LocalMux I__5813 (
            .O(N__27351),
            .I(N__27340));
    Span4Mux_h I__5812 (
            .O(N__27348),
            .I(N__27340));
    LocalMux I__5811 (
            .O(N__27345),
            .I(N__27337));
    Odrv4 I__5810 (
            .O(N__27340),
            .I(divider_4));
    Odrv12 I__5809 (
            .O(N__27337),
            .I(divider_4));
    InMux I__5808 (
            .O(N__27332),
            .I(N__27329));
    LocalMux I__5807 (
            .O(N__27329),
            .I(\Inst_core.Inst_sampler.n30 ));
    InMux I__5806 (
            .O(N__27326),
            .I(N__27323));
    LocalMux I__5805 (
            .O(N__27323),
            .I(N__27320));
    Odrv4 I__5804 (
            .O(N__27320),
            .I(\Inst_core.Inst_sampler.n8592 ));
    InMux I__5803 (
            .O(N__27317),
            .I(N__27310));
    InMux I__5802 (
            .O(N__27316),
            .I(N__27310));
    InMux I__5801 (
            .O(N__27315),
            .I(N__27307));
    LocalMux I__5800 (
            .O(N__27310),
            .I(N__27304));
    LocalMux I__5799 (
            .O(N__27307),
            .I(divider_2));
    Odrv12 I__5798 (
            .O(N__27304),
            .I(divider_2));
    InMux I__5797 (
            .O(N__27299),
            .I(N__27296));
    LocalMux I__5796 (
            .O(N__27296),
            .I(N__27291));
    InMux I__5795 (
            .O(N__27295),
            .I(N__27288));
    InMux I__5794 (
            .O(N__27294),
            .I(N__27285));
    Sp12to4 I__5793 (
            .O(N__27291),
            .I(N__27280));
    LocalMux I__5792 (
            .O(N__27288),
            .I(N__27280));
    LocalMux I__5791 (
            .O(N__27285),
            .I(divider_10));
    Odrv12 I__5790 (
            .O(N__27280),
            .I(divider_10));
    CascadeMux I__5789 (
            .O(N__27275),
            .I(N__27271));
    InMux I__5788 (
            .O(N__27274),
            .I(N__27266));
    InMux I__5787 (
            .O(N__27271),
            .I(N__27266));
    LocalMux I__5786 (
            .O(N__27266),
            .I(N__27263));
    Span4Mux_h I__5785 (
            .O(N__27263),
            .I(N__27259));
    InMux I__5784 (
            .O(N__27262),
            .I(N__27256));
    Span4Mux_v I__5783 (
            .O(N__27259),
            .I(N__27253));
    LocalMux I__5782 (
            .O(N__27256),
            .I(divider_8));
    Odrv4 I__5781 (
            .O(N__27253),
            .I(divider_8));
    CascadeMux I__5780 (
            .O(N__27248),
            .I(N__27244));
    InMux I__5779 (
            .O(N__27247),
            .I(N__27241));
    InMux I__5778 (
            .O(N__27244),
            .I(N__27238));
    LocalMux I__5777 (
            .O(N__27241),
            .I(N__27234));
    LocalMux I__5776 (
            .O(N__27238),
            .I(N__27231));
    InMux I__5775 (
            .O(N__27237),
            .I(N__27228));
    Span4Mux_v I__5774 (
            .O(N__27234),
            .I(N__27225));
    Span12Mux_s6_v I__5773 (
            .O(N__27231),
            .I(N__27222));
    LocalMux I__5772 (
            .O(N__27228),
            .I(divider_17));
    Odrv4 I__5771 (
            .O(N__27225),
            .I(divider_17));
    Odrv12 I__5770 (
            .O(N__27222),
            .I(divider_17));
    InMux I__5769 (
            .O(N__27215),
            .I(N__27212));
    LocalMux I__5768 (
            .O(N__27212),
            .I(\Inst_core.Inst_sampler.n8588 ));
    InMux I__5767 (
            .O(N__27209),
            .I(N__27202));
    CascadeMux I__5766 (
            .O(N__27208),
            .I(N__27194));
    InMux I__5765 (
            .O(N__27207),
            .I(N__27188));
    InMux I__5764 (
            .O(N__27206),
            .I(N__27183));
    InMux I__5763 (
            .O(N__27205),
            .I(N__27183));
    LocalMux I__5762 (
            .O(N__27202),
            .I(N__27180));
    InMux I__5761 (
            .O(N__27201),
            .I(N__27175));
    InMux I__5760 (
            .O(N__27200),
            .I(N__27175));
    InMux I__5759 (
            .O(N__27199),
            .I(N__27171));
    InMux I__5758 (
            .O(N__27198),
            .I(N__27168));
    InMux I__5757 (
            .O(N__27197),
            .I(N__27165));
    InMux I__5756 (
            .O(N__27194),
            .I(N__27162));
    InMux I__5755 (
            .O(N__27193),
            .I(N__27159));
    InMux I__5754 (
            .O(N__27192),
            .I(N__27156));
    InMux I__5753 (
            .O(N__27191),
            .I(N__27153));
    LocalMux I__5752 (
            .O(N__27188),
            .I(N__27150));
    LocalMux I__5751 (
            .O(N__27183),
            .I(N__27143));
    Span4Mux_s3_v I__5750 (
            .O(N__27180),
            .I(N__27143));
    LocalMux I__5749 (
            .O(N__27175),
            .I(N__27143));
    InMux I__5748 (
            .O(N__27174),
            .I(N__27137));
    LocalMux I__5747 (
            .O(N__27171),
            .I(N__27134));
    LocalMux I__5746 (
            .O(N__27168),
            .I(N__27129));
    LocalMux I__5745 (
            .O(N__27165),
            .I(N__27129));
    LocalMux I__5744 (
            .O(N__27162),
            .I(N__27124));
    LocalMux I__5743 (
            .O(N__27159),
            .I(N__27124));
    LocalMux I__5742 (
            .O(N__27156),
            .I(N__27121));
    LocalMux I__5741 (
            .O(N__27153),
            .I(N__27114));
    Span4Mux_v I__5740 (
            .O(N__27150),
            .I(N__27114));
    Span4Mux_v I__5739 (
            .O(N__27143),
            .I(N__27114));
    InMux I__5738 (
            .O(N__27142),
            .I(N__27107));
    InMux I__5737 (
            .O(N__27141),
            .I(N__27107));
    InMux I__5736 (
            .O(N__27140),
            .I(N__27107));
    LocalMux I__5735 (
            .O(N__27137),
            .I(N__27104));
    Span4Mux_v I__5734 (
            .O(N__27134),
            .I(N__27101));
    Span4Mux_h I__5733 (
            .O(N__27129),
            .I(N__27098));
    Span4Mux_h I__5732 (
            .O(N__27124),
            .I(N__27095));
    Span4Mux_h I__5731 (
            .O(N__27121),
            .I(N__27090));
    Span4Mux_h I__5730 (
            .O(N__27114),
            .I(N__27090));
    LocalMux I__5729 (
            .O(N__27107),
            .I(cmd_15));
    Odrv4 I__5728 (
            .O(N__27104),
            .I(cmd_15));
    Odrv4 I__5727 (
            .O(N__27101),
            .I(cmd_15));
    Odrv4 I__5726 (
            .O(N__27098),
            .I(cmd_15));
    Odrv4 I__5725 (
            .O(N__27095),
            .I(cmd_15));
    Odrv4 I__5724 (
            .O(N__27090),
            .I(cmd_15));
    InMux I__5723 (
            .O(N__27077),
            .I(N__27073));
    InMux I__5722 (
            .O(N__27076),
            .I(N__27070));
    LocalMux I__5721 (
            .O(N__27073),
            .I(bwd_7));
    LocalMux I__5720 (
            .O(N__27070),
            .I(bwd_7));
    InMux I__5719 (
            .O(N__27065),
            .I(N__27061));
    InMux I__5718 (
            .O(N__27064),
            .I(N__27058));
    LocalMux I__5717 (
            .O(N__27061),
            .I(fwd_10));
    LocalMux I__5716 (
            .O(N__27058),
            .I(fwd_10));
    InMux I__5715 (
            .O(N__27053),
            .I(N__27044));
    InMux I__5714 (
            .O(N__27052),
            .I(N__27044));
    InMux I__5713 (
            .O(N__27051),
            .I(N__27039));
    InMux I__5712 (
            .O(N__27050),
            .I(N__27036));
    InMux I__5711 (
            .O(N__27049),
            .I(N__27033));
    LocalMux I__5710 (
            .O(N__27044),
            .I(N__27030));
    InMux I__5709 (
            .O(N__27043),
            .I(N__27027));
    InMux I__5708 (
            .O(N__27042),
            .I(N__27024));
    LocalMux I__5707 (
            .O(N__27039),
            .I(N__27018));
    LocalMux I__5706 (
            .O(N__27036),
            .I(N__27018));
    LocalMux I__5705 (
            .O(N__27033),
            .I(N__27015));
    Span4Mux_v I__5704 (
            .O(N__27030),
            .I(N__27008));
    LocalMux I__5703 (
            .O(N__27027),
            .I(N__27008));
    LocalMux I__5702 (
            .O(N__27024),
            .I(N__27008));
    InMux I__5701 (
            .O(N__27023),
            .I(N__27005));
    Span4Mux_h I__5700 (
            .O(N__27018),
            .I(N__27002));
    Span4Mux_s3_h I__5699 (
            .O(N__27015),
            .I(N__26997));
    Span4Mux_v I__5698 (
            .O(N__27008),
            .I(N__26997));
    LocalMux I__5697 (
            .O(N__27005),
            .I(N__26994));
    Span4Mux_v I__5696 (
            .O(N__27002),
            .I(N__26991));
    Span4Mux_h I__5695 (
            .O(N__26997),
            .I(N__26988));
    Odrv4 I__5694 (
            .O(N__26994),
            .I(wrtrigmask_2));
    Odrv4 I__5693 (
            .O(N__26991),
            .I(wrtrigmask_2));
    Odrv4 I__5692 (
            .O(N__26988),
            .I(wrtrigmask_2));
    InMux I__5691 (
            .O(N__26981),
            .I(N__26977));
    InMux I__5690 (
            .O(N__26980),
            .I(N__26974));
    LocalMux I__5689 (
            .O(N__26977),
            .I(maskRegister_4_adj_1324));
    LocalMux I__5688 (
            .O(N__26974),
            .I(maskRegister_4_adj_1324));
    CascadeMux I__5687 (
            .O(N__26969),
            .I(N__26966));
    InMux I__5686 (
            .O(N__26966),
            .I(N__26963));
    LocalMux I__5685 (
            .O(N__26963),
            .I(N__26959));
    InMux I__5684 (
            .O(N__26962),
            .I(N__26956));
    Span4Mux_h I__5683 (
            .O(N__26959),
            .I(N__26953));
    LocalMux I__5682 (
            .O(N__26956),
            .I(\Inst_core.Inst_sync.filteredInput_7 ));
    Odrv4 I__5681 (
            .O(N__26953),
            .I(\Inst_core.Inst_sync.filteredInput_7 ));
    SRMux I__5680 (
            .O(N__26948),
            .I(N__26945));
    LocalMux I__5679 (
            .O(N__26945),
            .I(N__26942));
    Span4Mux_h I__5678 (
            .O(N__26942),
            .I(N__26939));
    Odrv4 I__5677 (
            .O(N__26939),
            .I(\Inst_core.Inst_sync.Inst_filter.n4735 ));
    InMux I__5676 (
            .O(N__26936),
            .I(N__26933));
    LocalMux I__5675 (
            .O(N__26933),
            .I(N__26929));
    InMux I__5674 (
            .O(N__26932),
            .I(N__26926));
    Span4Mux_h I__5673 (
            .O(N__26929),
            .I(N__26923));
    LocalMux I__5672 (
            .O(N__26926),
            .I(maskRegister_7_adj_1281));
    Odrv4 I__5671 (
            .O(N__26923),
            .I(maskRegister_7_adj_1281));
    SRMux I__5670 (
            .O(N__26918),
            .I(N__26915));
    LocalMux I__5669 (
            .O(N__26915),
            .I(N__26912));
    Sp12to4 I__5668 (
            .O(N__26912),
            .I(N__26909));
    Span12Mux_s0_v I__5667 (
            .O(N__26909),
            .I(N__26906));
    Odrv12 I__5666 (
            .O(N__26906),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4752 ));
    InMux I__5665 (
            .O(N__26903),
            .I(N__26899));
    InMux I__5664 (
            .O(N__26902),
            .I(N__26896));
    LocalMux I__5663 (
            .O(N__26899),
            .I(N__26893));
    LocalMux I__5662 (
            .O(N__26896),
            .I(maskRegister_0_adj_1328));
    Odrv4 I__5661 (
            .O(N__26893),
            .I(maskRegister_0_adj_1328));
    InMux I__5660 (
            .O(N__26888),
            .I(N__26884));
    InMux I__5659 (
            .O(N__26887),
            .I(N__26881));
    LocalMux I__5658 (
            .O(N__26884),
            .I(N__26878));
    LocalMux I__5657 (
            .O(N__26881),
            .I(bwd_9));
    Odrv4 I__5656 (
            .O(N__26878),
            .I(bwd_9));
    InMux I__5655 (
            .O(N__26873),
            .I(N__26870));
    LocalMux I__5654 (
            .O(N__26870),
            .I(\Inst_core.Inst_controller.n24 ));
    CascadeMux I__5653 (
            .O(N__26867),
            .I(\Inst_core.Inst_controller.n22_adj_988_cascade_ ));
    InMux I__5652 (
            .O(N__26864),
            .I(N__26861));
    LocalMux I__5651 (
            .O(N__26861),
            .I(N__26858));
    Span4Mux_h I__5650 (
            .O(N__26858),
            .I(N__26853));
    InMux I__5649 (
            .O(N__26857),
            .I(N__26848));
    InMux I__5648 (
            .O(N__26856),
            .I(N__26848));
    Odrv4 I__5647 (
            .O(N__26853),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3 ));
    LocalMux I__5646 (
            .O(N__26848),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3 ));
    InMux I__5645 (
            .O(N__26843),
            .I(N__26839));
    InMux I__5644 (
            .O(N__26842),
            .I(N__26836));
    LocalMux I__5643 (
            .O(N__26839),
            .I(valueRegister_3_adj_1293));
    LocalMux I__5642 (
            .O(N__26836),
            .I(valueRegister_3_adj_1293));
    CascadeMux I__5641 (
            .O(N__26831),
            .I(N__26828));
    InMux I__5640 (
            .O(N__26828),
            .I(N__26825));
    LocalMux I__5639 (
            .O(N__26825),
            .I(N__26822));
    Span4Mux_h I__5638 (
            .O(N__26822),
            .I(N__26819));
    Span4Mux_h I__5637 (
            .O(N__26819),
            .I(N__26816));
    Odrv4 I__5636 (
            .O(N__26816),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_3 ));
    SRMux I__5635 (
            .O(N__26813),
            .I(N__26810));
    LocalMux I__5634 (
            .O(N__26810),
            .I(N__26807));
    Span4Mux_h I__5633 (
            .O(N__26807),
            .I(N__26804));
    Odrv4 I__5632 (
            .O(N__26804),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4748 ));
    InMux I__5631 (
            .O(N__26801),
            .I(N__26797));
    InMux I__5630 (
            .O(N__26800),
            .I(N__26794));
    LocalMux I__5629 (
            .O(N__26797),
            .I(bwd_6));
    LocalMux I__5628 (
            .O(N__26794),
            .I(bwd_6));
    CascadeMux I__5627 (
            .O(N__26789),
            .I(N__26786));
    InMux I__5626 (
            .O(N__26786),
            .I(N__26782));
    InMux I__5625 (
            .O(N__26785),
            .I(N__26779));
    LocalMux I__5624 (
            .O(N__26782),
            .I(N__26776));
    LocalMux I__5623 (
            .O(N__26779),
            .I(bwd_5));
    Odrv4 I__5622 (
            .O(N__26776),
            .I(bwd_5));
    InMux I__5621 (
            .O(N__26771),
            .I(N__26768));
    LocalMux I__5620 (
            .O(N__26768),
            .I(\Inst_core.Inst_controller.n23 ));
    InMux I__5619 (
            .O(N__26765),
            .I(N__26761));
    InMux I__5618 (
            .O(N__26764),
            .I(N__26758));
    LocalMux I__5617 (
            .O(N__26761),
            .I(bwd_3));
    LocalMux I__5616 (
            .O(N__26758),
            .I(bwd_3));
    CascadeMux I__5615 (
            .O(N__26753),
            .I(N__26749));
    InMux I__5614 (
            .O(N__26752),
            .I(N__26746));
    InMux I__5613 (
            .O(N__26749),
            .I(N__26743));
    LocalMux I__5612 (
            .O(N__26746),
            .I(bwd_4));
    LocalMux I__5611 (
            .O(N__26743),
            .I(bwd_4));
    InMux I__5610 (
            .O(N__26738),
            .I(N__26735));
    LocalMux I__5609 (
            .O(N__26735),
            .I(\Inst_core.Inst_controller.n21_adj_989 ));
    CascadeMux I__5608 (
            .O(N__26732),
            .I(N__26722));
    InMux I__5607 (
            .O(N__26731),
            .I(N__26717));
    InMux I__5606 (
            .O(N__26730),
            .I(N__26713));
    InMux I__5605 (
            .O(N__26729),
            .I(N__26702));
    InMux I__5604 (
            .O(N__26728),
            .I(N__26702));
    InMux I__5603 (
            .O(N__26727),
            .I(N__26702));
    InMux I__5602 (
            .O(N__26726),
            .I(N__26702));
    InMux I__5601 (
            .O(N__26725),
            .I(N__26699));
    InMux I__5600 (
            .O(N__26722),
            .I(N__26691));
    InMux I__5599 (
            .O(N__26721),
            .I(N__26691));
    InMux I__5598 (
            .O(N__26720),
            .I(N__26691));
    LocalMux I__5597 (
            .O(N__26717),
            .I(N__26688));
    InMux I__5596 (
            .O(N__26716),
            .I(N__26685));
    LocalMux I__5595 (
            .O(N__26713),
            .I(N__26682));
    InMux I__5594 (
            .O(N__26712),
            .I(N__26677));
    InMux I__5593 (
            .O(N__26711),
            .I(N__26677));
    LocalMux I__5592 (
            .O(N__26702),
            .I(N__26674));
    LocalMux I__5591 (
            .O(N__26699),
            .I(N__26671));
    InMux I__5590 (
            .O(N__26698),
            .I(N__26668));
    LocalMux I__5589 (
            .O(N__26691),
            .I(N__26665));
    Span4Mux_h I__5588 (
            .O(N__26688),
            .I(N__26660));
    LocalMux I__5587 (
            .O(N__26685),
            .I(N__26660));
    Span4Mux_v I__5586 (
            .O(N__26682),
            .I(N__26655));
    LocalMux I__5585 (
            .O(N__26677),
            .I(N__26655));
    Span4Mux_v I__5584 (
            .O(N__26674),
            .I(N__26649));
    Span4Mux_h I__5583 (
            .O(N__26671),
            .I(N__26646));
    LocalMux I__5582 (
            .O(N__26668),
            .I(N__26643));
    Span4Mux_s2_v I__5581 (
            .O(N__26665),
            .I(N__26636));
    Span4Mux_v I__5580 (
            .O(N__26660),
            .I(N__26636));
    Span4Mux_h I__5579 (
            .O(N__26655),
            .I(N__26636));
    InMux I__5578 (
            .O(N__26654),
            .I(N__26633));
    InMux I__5577 (
            .O(N__26653),
            .I(N__26630));
    InMux I__5576 (
            .O(N__26652),
            .I(N__26627));
    Odrv4 I__5575 (
            .O(N__26649),
            .I(cmd_11));
    Odrv4 I__5574 (
            .O(N__26646),
            .I(cmd_11));
    Odrv4 I__5573 (
            .O(N__26643),
            .I(cmd_11));
    Odrv4 I__5572 (
            .O(N__26636),
            .I(cmd_11));
    LocalMux I__5571 (
            .O(N__26633),
            .I(cmd_11));
    LocalMux I__5570 (
            .O(N__26630),
            .I(cmd_11));
    LocalMux I__5569 (
            .O(N__26627),
            .I(cmd_11));
    InMux I__5568 (
            .O(N__26612),
            .I(N__26608));
    InMux I__5567 (
            .O(N__26611),
            .I(N__26605));
    LocalMux I__5566 (
            .O(N__26608),
            .I(N__26602));
    LocalMux I__5565 (
            .O(N__26605),
            .I(configRegister_16_adj_1304));
    Odrv4 I__5564 (
            .O(N__26602),
            .I(configRegister_16_adj_1304));
    InMux I__5563 (
            .O(N__26597),
            .I(N__26591));
    InMux I__5562 (
            .O(N__26596),
            .I(N__26588));
    InMux I__5561 (
            .O(N__26595),
            .I(N__26579));
    InMux I__5560 (
            .O(N__26594),
            .I(N__26579));
    LocalMux I__5559 (
            .O(N__26591),
            .I(N__26576));
    LocalMux I__5558 (
            .O(N__26588),
            .I(N__26573));
    InMux I__5557 (
            .O(N__26587),
            .I(N__26570));
    InMux I__5556 (
            .O(N__26586),
            .I(N__26567));
    InMux I__5555 (
            .O(N__26585),
            .I(N__26564));
    InMux I__5554 (
            .O(N__26584),
            .I(N__26561));
    LocalMux I__5553 (
            .O(N__26579),
            .I(N__26556));
    Span4Mux_h I__5552 (
            .O(N__26576),
            .I(N__26556));
    Span4Mux_v I__5551 (
            .O(N__26573),
            .I(N__26553));
    LocalMux I__5550 (
            .O(N__26570),
            .I(cmd_17));
    LocalMux I__5549 (
            .O(N__26567),
            .I(cmd_17));
    LocalMux I__5548 (
            .O(N__26564),
            .I(cmd_17));
    LocalMux I__5547 (
            .O(N__26561),
            .I(cmd_17));
    Odrv4 I__5546 (
            .O(N__26556),
            .I(cmd_17));
    Odrv4 I__5545 (
            .O(N__26553),
            .I(cmd_17));
    InMux I__5544 (
            .O(N__26540),
            .I(N__26537));
    LocalMux I__5543 (
            .O(N__26537),
            .I(N__26531));
    InMux I__5542 (
            .O(N__26536),
            .I(N__26528));
    InMux I__5541 (
            .O(N__26535),
            .I(N__26525));
    CascadeMux I__5540 (
            .O(N__26534),
            .I(N__26521));
    Span4Mux_h I__5539 (
            .O(N__26531),
            .I(N__26515));
    LocalMux I__5538 (
            .O(N__26528),
            .I(N__26512));
    LocalMux I__5537 (
            .O(N__26525),
            .I(N__26509));
    InMux I__5536 (
            .O(N__26524),
            .I(N__26504));
    InMux I__5535 (
            .O(N__26521),
            .I(N__26504));
    InMux I__5534 (
            .O(N__26520),
            .I(N__26497));
    InMux I__5533 (
            .O(N__26519),
            .I(N__26497));
    InMux I__5532 (
            .O(N__26518),
            .I(N__26497));
    Odrv4 I__5531 (
            .O(N__26515),
            .I(cmd_28));
    Odrv4 I__5530 (
            .O(N__26512),
            .I(cmd_28));
    Odrv4 I__5529 (
            .O(N__26509),
            .I(cmd_28));
    LocalMux I__5528 (
            .O(N__26504),
            .I(cmd_28));
    LocalMux I__5527 (
            .O(N__26497),
            .I(cmd_28));
    CascadeMux I__5526 (
            .O(N__26486),
            .I(N__26482));
    InMux I__5525 (
            .O(N__26485),
            .I(N__26479));
    InMux I__5524 (
            .O(N__26482),
            .I(N__26476));
    LocalMux I__5523 (
            .O(N__26479),
            .I(fwd_3));
    LocalMux I__5522 (
            .O(N__26476),
            .I(fwd_3));
    InMux I__5521 (
            .O(N__26471),
            .I(N__26467));
    InMux I__5520 (
            .O(N__26470),
            .I(N__26464));
    LocalMux I__5519 (
            .O(N__26467),
            .I(N__26461));
    LocalMux I__5518 (
            .O(N__26464),
            .I(maskRegister_7_adj_1321));
    Odrv12 I__5517 (
            .O(N__26461),
            .I(maskRegister_7_adj_1321));
    SRMux I__5516 (
            .O(N__26456),
            .I(N__26453));
    LocalMux I__5515 (
            .O(N__26453),
            .I(N__26450));
    Span4Mux_h I__5514 (
            .O(N__26450),
            .I(N__26447));
    Span4Mux_v I__5513 (
            .O(N__26447),
            .I(N__26444));
    Odrv4 I__5512 (
            .O(N__26444),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4759 ));
    InMux I__5511 (
            .O(N__26441),
            .I(N__26438));
    LocalMux I__5510 (
            .O(N__26438),
            .I(N__26434));
    InMux I__5509 (
            .O(N__26437),
            .I(N__26431));
    Odrv4 I__5508 (
            .O(N__26434),
            .I(maskRegister_0_adj_1368));
    LocalMux I__5507 (
            .O(N__26431),
            .I(maskRegister_0_adj_1368));
    InMux I__5506 (
            .O(N__26426),
            .I(N__26422));
    InMux I__5505 (
            .O(N__26425),
            .I(N__26419));
    LocalMux I__5504 (
            .O(N__26422),
            .I(maskRegister_1_adj_1367));
    LocalMux I__5503 (
            .O(N__26419),
            .I(maskRegister_1_adj_1367));
    InMux I__5502 (
            .O(N__26414),
            .I(N__26410));
    InMux I__5501 (
            .O(N__26413),
            .I(N__26407));
    LocalMux I__5500 (
            .O(N__26410),
            .I(maskRegister_2_adj_1366));
    LocalMux I__5499 (
            .O(N__26407),
            .I(maskRegister_2_adj_1366));
    InMux I__5498 (
            .O(N__26402),
            .I(N__26399));
    LocalMux I__5497 (
            .O(N__26399),
            .I(N__26396));
    Span4Mux_v I__5496 (
            .O(N__26396),
            .I(N__26393));
    Odrv4 I__5495 (
            .O(N__26393),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7_adj_996 ));
    InMux I__5494 (
            .O(N__26390),
            .I(N__26363));
    InMux I__5493 (
            .O(N__26389),
            .I(N__26363));
    InMux I__5492 (
            .O(N__26388),
            .I(N__26363));
    InMux I__5491 (
            .O(N__26387),
            .I(N__26363));
    InMux I__5490 (
            .O(N__26386),
            .I(N__26363));
    InMux I__5489 (
            .O(N__26385),
            .I(N__26363));
    InMux I__5488 (
            .O(N__26384),
            .I(N__26363));
    InMux I__5487 (
            .O(N__26383),
            .I(N__26363));
    InMux I__5486 (
            .O(N__26382),
            .I(N__26346));
    InMux I__5485 (
            .O(N__26381),
            .I(N__26343));
    InMux I__5484 (
            .O(N__26380),
            .I(N__26332));
    LocalMux I__5483 (
            .O(N__26363),
            .I(N__26329));
    InMux I__5482 (
            .O(N__26362),
            .I(N__26326));
    InMux I__5481 (
            .O(N__26361),
            .I(N__26315));
    InMux I__5480 (
            .O(N__26360),
            .I(N__26315));
    InMux I__5479 (
            .O(N__26359),
            .I(N__26315));
    InMux I__5478 (
            .O(N__26358),
            .I(N__26315));
    InMux I__5477 (
            .O(N__26357),
            .I(N__26315));
    InMux I__5476 (
            .O(N__26356),
            .I(N__26298));
    InMux I__5475 (
            .O(N__26355),
            .I(N__26298));
    InMux I__5474 (
            .O(N__26354),
            .I(N__26298));
    InMux I__5473 (
            .O(N__26353),
            .I(N__26298));
    InMux I__5472 (
            .O(N__26352),
            .I(N__26298));
    InMux I__5471 (
            .O(N__26351),
            .I(N__26298));
    InMux I__5470 (
            .O(N__26350),
            .I(N__26298));
    InMux I__5469 (
            .O(N__26349),
            .I(N__26298));
    LocalMux I__5468 (
            .O(N__26346),
            .I(N__26295));
    LocalMux I__5467 (
            .O(N__26343),
            .I(N__26292));
    InMux I__5466 (
            .O(N__26342),
            .I(N__26274));
    InMux I__5465 (
            .O(N__26341),
            .I(N__26274));
    InMux I__5464 (
            .O(N__26340),
            .I(N__26274));
    InMux I__5463 (
            .O(N__26339),
            .I(N__26274));
    InMux I__5462 (
            .O(N__26338),
            .I(N__26274));
    InMux I__5461 (
            .O(N__26337),
            .I(N__26274));
    InMux I__5460 (
            .O(N__26336),
            .I(N__26274));
    InMux I__5459 (
            .O(N__26335),
            .I(N__26274));
    LocalMux I__5458 (
            .O(N__26332),
            .I(N__26271));
    Span4Mux_s2_v I__5457 (
            .O(N__26329),
            .I(N__26256));
    LocalMux I__5456 (
            .O(N__26326),
            .I(N__26256));
    LocalMux I__5455 (
            .O(N__26315),
            .I(N__26256));
    LocalMux I__5454 (
            .O(N__26298),
            .I(N__26253));
    Span4Mux_v I__5453 (
            .O(N__26295),
            .I(N__26248));
    Span4Mux_v I__5452 (
            .O(N__26292),
            .I(N__26248));
    InMux I__5451 (
            .O(N__26291),
            .I(N__26245));
    LocalMux I__5450 (
            .O(N__26274),
            .I(N__26241));
    Span4Mux_h I__5449 (
            .O(N__26271),
            .I(N__26238));
    InMux I__5448 (
            .O(N__26270),
            .I(N__26221));
    InMux I__5447 (
            .O(N__26269),
            .I(N__26221));
    InMux I__5446 (
            .O(N__26268),
            .I(N__26221));
    InMux I__5445 (
            .O(N__26267),
            .I(N__26221));
    InMux I__5444 (
            .O(N__26266),
            .I(N__26221));
    InMux I__5443 (
            .O(N__26265),
            .I(N__26221));
    InMux I__5442 (
            .O(N__26264),
            .I(N__26221));
    InMux I__5441 (
            .O(N__26263),
            .I(N__26221));
    Span4Mux_v I__5440 (
            .O(N__26256),
            .I(N__26218));
    Span4Mux_v I__5439 (
            .O(N__26253),
            .I(N__26211));
    Span4Mux_h I__5438 (
            .O(N__26248),
            .I(N__26211));
    LocalMux I__5437 (
            .O(N__26245),
            .I(N__26211));
    InMux I__5436 (
            .O(N__26244),
            .I(N__26208));
    Span4Mux_h I__5435 (
            .O(N__26241),
            .I(N__26203));
    Span4Mux_v I__5434 (
            .O(N__26238),
            .I(N__26203));
    LocalMux I__5433 (
            .O(N__26221),
            .I(N__26198));
    Span4Mux_h I__5432 (
            .O(N__26218),
            .I(N__26198));
    Odrv4 I__5431 (
            .O(N__26211),
            .I(flagDemux));
    LocalMux I__5430 (
            .O(N__26208),
            .I(flagDemux));
    Odrv4 I__5429 (
            .O(N__26203),
            .I(flagDemux));
    Odrv4 I__5428 (
            .O(N__26198),
            .I(flagDemux));
    InMux I__5427 (
            .O(N__26189),
            .I(N__26183));
    InMux I__5426 (
            .O(N__26188),
            .I(N__26183));
    LocalMux I__5425 (
            .O(N__26183),
            .I(N__26180));
    Odrv12 I__5424 (
            .O(N__26180),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register ));
    InMux I__5423 (
            .O(N__26177),
            .I(N__26174));
    LocalMux I__5422 (
            .O(N__26174),
            .I(N__26170));
    InMux I__5421 (
            .O(N__26173),
            .I(N__26167));
    Odrv4 I__5420 (
            .O(N__26170),
            .I(valueRegister_5_adj_1371));
    LocalMux I__5419 (
            .O(N__26167),
            .I(valueRegister_5_adj_1371));
    InMux I__5418 (
            .O(N__26162),
            .I(N__26159));
    LocalMux I__5417 (
            .O(N__26159),
            .I(N__26156));
    Span4Mux_h I__5416 (
            .O(N__26156),
            .I(N__26152));
    InMux I__5415 (
            .O(N__26155),
            .I(N__26149));
    Odrv4 I__5414 (
            .O(N__26152),
            .I(configRegister_13_adj_1387));
    LocalMux I__5413 (
            .O(N__26149),
            .I(configRegister_13_adj_1387));
    InMux I__5412 (
            .O(N__26144),
            .I(N__26138));
    InMux I__5411 (
            .O(N__26143),
            .I(N__26138));
    LocalMux I__5410 (
            .O(N__26138),
            .I(N__26131));
    InMux I__5409 (
            .O(N__26137),
            .I(N__26128));
    InMux I__5408 (
            .O(N__26136),
            .I(N__26124));
    CascadeMux I__5407 (
            .O(N__26135),
            .I(N__26121));
    CascadeMux I__5406 (
            .O(N__26134),
            .I(N__26115));
    Span4Mux_v I__5405 (
            .O(N__26131),
            .I(N__26107));
    LocalMux I__5404 (
            .O(N__26128),
            .I(N__26107));
    InMux I__5403 (
            .O(N__26127),
            .I(N__26103));
    LocalMux I__5402 (
            .O(N__26124),
            .I(N__26097));
    InMux I__5401 (
            .O(N__26121),
            .I(N__26092));
    InMux I__5400 (
            .O(N__26120),
            .I(N__26092));
    InMux I__5399 (
            .O(N__26119),
            .I(N__26089));
    InMux I__5398 (
            .O(N__26118),
            .I(N__26077));
    InMux I__5397 (
            .O(N__26115),
            .I(N__26077));
    InMux I__5396 (
            .O(N__26114),
            .I(N__26077));
    InMux I__5395 (
            .O(N__26113),
            .I(N__26077));
    InMux I__5394 (
            .O(N__26112),
            .I(N__26072));
    Span4Mux_v I__5393 (
            .O(N__26107),
            .I(N__26069));
    InMux I__5392 (
            .O(N__26106),
            .I(N__26066));
    LocalMux I__5391 (
            .O(N__26103),
            .I(N__26063));
    InMux I__5390 (
            .O(N__26102),
            .I(N__26060));
    InMux I__5389 (
            .O(N__26101),
            .I(N__26055));
    InMux I__5388 (
            .O(N__26100),
            .I(N__26055));
    Span4Mux_v I__5387 (
            .O(N__26097),
            .I(N__26050));
    LocalMux I__5386 (
            .O(N__26092),
            .I(N__26050));
    LocalMux I__5385 (
            .O(N__26089),
            .I(N__26045));
    InMux I__5384 (
            .O(N__26088),
            .I(N__26038));
    InMux I__5383 (
            .O(N__26087),
            .I(N__26038));
    InMux I__5382 (
            .O(N__26086),
            .I(N__26038));
    LocalMux I__5381 (
            .O(N__26077),
            .I(N__26035));
    InMux I__5380 (
            .O(N__26076),
            .I(N__26030));
    InMux I__5379 (
            .O(N__26075),
            .I(N__26030));
    LocalMux I__5378 (
            .O(N__26072),
            .I(N__26027));
    Sp12to4 I__5377 (
            .O(N__26069),
            .I(N__26021));
    LocalMux I__5376 (
            .O(N__26066),
            .I(N__26021));
    Span4Mux_v I__5375 (
            .O(N__26063),
            .I(N__26012));
    LocalMux I__5374 (
            .O(N__26060),
            .I(N__26012));
    LocalMux I__5373 (
            .O(N__26055),
            .I(N__26012));
    Span4Mux_h I__5372 (
            .O(N__26050),
            .I(N__26012));
    InMux I__5371 (
            .O(N__26049),
            .I(N__26007));
    InMux I__5370 (
            .O(N__26048),
            .I(N__26007));
    Span4Mux_v I__5369 (
            .O(N__26045),
            .I(N__26000));
    LocalMux I__5368 (
            .O(N__26038),
            .I(N__26000));
    Span4Mux_s1_v I__5367 (
            .O(N__26035),
            .I(N__26000));
    LocalMux I__5366 (
            .O(N__26030),
            .I(N__25995));
    Span4Mux_v I__5365 (
            .O(N__26027),
            .I(N__25995));
    InMux I__5364 (
            .O(N__26026),
            .I(N__25992));
    Span12Mux_s8_h I__5363 (
            .O(N__26021),
            .I(N__25989));
    Span4Mux_h I__5362 (
            .O(N__26012),
            .I(N__25986));
    LocalMux I__5361 (
            .O(N__26007),
            .I(N__25979));
    Span4Mux_v I__5360 (
            .O(N__26000),
            .I(N__25979));
    Span4Mux_h I__5359 (
            .O(N__25995),
            .I(N__25979));
    LocalMux I__5358 (
            .O(N__25992),
            .I(wrtrigcfg_3));
    Odrv12 I__5357 (
            .O(N__25989),
            .I(wrtrigcfg_3));
    Odrv4 I__5356 (
            .O(N__25986),
            .I(wrtrigcfg_3));
    Odrv4 I__5355 (
            .O(N__25979),
            .I(wrtrigcfg_3));
    InMux I__5354 (
            .O(N__25970),
            .I(N__25966));
    InMux I__5353 (
            .O(N__25969),
            .I(N__25963));
    LocalMux I__5352 (
            .O(N__25966),
            .I(N__25960));
    LocalMux I__5351 (
            .O(N__25963),
            .I(configRegister_16_adj_1384));
    Odrv4 I__5350 (
            .O(N__25960),
            .I(configRegister_16_adj_1384));
    InMux I__5349 (
            .O(N__25955),
            .I(N__25952));
    LocalMux I__5348 (
            .O(N__25952),
            .I(N__25948));
    InMux I__5347 (
            .O(N__25951),
            .I(N__25945));
    Odrv4 I__5346 (
            .O(N__25948),
            .I(configRegister_12_adj_1348));
    LocalMux I__5345 (
            .O(N__25945),
            .I(configRegister_12_adj_1348));
    SRMux I__5344 (
            .O(N__25940),
            .I(N__25929));
    InMux I__5343 (
            .O(N__25939),
            .I(N__25920));
    InMux I__5342 (
            .O(N__25938),
            .I(N__25920));
    InMux I__5341 (
            .O(N__25937),
            .I(N__25920));
    InMux I__5340 (
            .O(N__25936),
            .I(N__25920));
    InMux I__5339 (
            .O(N__25935),
            .I(N__25911));
    InMux I__5338 (
            .O(N__25934),
            .I(N__25911));
    InMux I__5337 (
            .O(N__25933),
            .I(N__25911));
    InMux I__5336 (
            .O(N__25932),
            .I(N__25911));
    LocalMux I__5335 (
            .O(N__25929),
            .I(N__25908));
    LocalMux I__5334 (
            .O(N__25920),
            .I(N__25903));
    LocalMux I__5333 (
            .O(N__25911),
            .I(N__25903));
    Span12Mux_s11_v I__5332 (
            .O(N__25908),
            .I(N__25898));
    Span12Mux_s4_v I__5331 (
            .O(N__25903),
            .I(N__25898));
    Odrv12 I__5330 (
            .O(N__25898),
            .I(\Inst_core.arm ));
    InMux I__5329 (
            .O(N__25895),
            .I(N__25891));
    InMux I__5328 (
            .O(N__25894),
            .I(N__25888));
    LocalMux I__5327 (
            .O(N__25891),
            .I(maskRegister_5_adj_1323));
    LocalMux I__5326 (
            .O(N__25888),
            .I(maskRegister_5_adj_1323));
    SRMux I__5325 (
            .O(N__25883),
            .I(N__25880));
    LocalMux I__5324 (
            .O(N__25880),
            .I(N__25877));
    Span4Mux_h I__5323 (
            .O(N__25877),
            .I(N__25874));
    Span4Mux_v I__5322 (
            .O(N__25874),
            .I(N__25871));
    Odrv4 I__5321 (
            .O(N__25871),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4757 ));
    InMux I__5320 (
            .O(N__25868),
            .I(N__25864));
    InMux I__5319 (
            .O(N__25867),
            .I(N__25861));
    LocalMux I__5318 (
            .O(N__25864),
            .I(maskRegister_6_adj_1322));
    LocalMux I__5317 (
            .O(N__25861),
            .I(maskRegister_6_adj_1322));
    CascadeMux I__5316 (
            .O(N__25856),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n2_cascade_ ));
    InMux I__5315 (
            .O(N__25853),
            .I(N__25850));
    LocalMux I__5314 (
            .O(N__25850),
            .I(N__25847));
    Span4Mux_v I__5313 (
            .O(N__25847),
            .I(N__25844));
    Odrv4 I__5312 (
            .O(N__25844),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register ));
    InMux I__5311 (
            .O(N__25841),
            .I(N__25838));
    LocalMux I__5310 (
            .O(N__25838),
            .I(N__25835));
    Odrv4 I__5309 (
            .O(N__25835),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n100 ));
    InMux I__5308 (
            .O(N__25832),
            .I(N__25828));
    InMux I__5307 (
            .O(N__25831),
            .I(N__25825));
    LocalMux I__5306 (
            .O(N__25828),
            .I(N__25822));
    LocalMux I__5305 (
            .O(N__25825),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n553 ));
    Odrv4 I__5304 (
            .O(N__25822),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n553 ));
    CascadeMux I__5303 (
            .O(N__25817),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n100_cascade_ ));
    InMux I__5302 (
            .O(N__25814),
            .I(N__25811));
    LocalMux I__5301 (
            .O(N__25811),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register ));
    CascadeMux I__5300 (
            .O(N__25808),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n2_cascade_ ));
    InMux I__5299 (
            .O(N__25805),
            .I(N__25802));
    LocalMux I__5298 (
            .O(N__25802),
            .I(N__25798));
    InMux I__5297 (
            .O(N__25801),
            .I(N__25795));
    Span4Mux_s3_h I__5296 (
            .O(N__25798),
            .I(N__25792));
    LocalMux I__5295 (
            .O(N__25795),
            .I(configRegister_17_adj_1383));
    Odrv4 I__5294 (
            .O(N__25792),
            .I(configRegister_17_adj_1383));
    InMux I__5293 (
            .O(N__25787),
            .I(N__25784));
    LocalMux I__5292 (
            .O(N__25784),
            .I(N__25781));
    Odrv4 I__5291 (
            .O(N__25781),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n100 ));
    CascadeMux I__5290 (
            .O(N__25778),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n100_cascade_ ));
    CascadeMux I__5289 (
            .O(N__25775),
            .I(N__25771));
    InMux I__5288 (
            .O(N__25774),
            .I(N__25768));
    InMux I__5287 (
            .O(N__25771),
            .I(N__25765));
    LocalMux I__5286 (
            .O(N__25768),
            .I(N__25762));
    LocalMux I__5285 (
            .O(N__25765),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n759 ));
    Odrv4 I__5284 (
            .O(N__25762),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n759 ));
    InMux I__5283 (
            .O(N__25757),
            .I(N__25754));
    LocalMux I__5282 (
            .O(N__25754),
            .I(N__25751));
    Odrv4 I__5281 (
            .O(N__25751),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n770 ));
    CascadeMux I__5280 (
            .O(N__25748),
            .I(N__25740));
    InMux I__5279 (
            .O(N__25747),
            .I(N__25736));
    InMux I__5278 (
            .O(N__25746),
            .I(N__25727));
    InMux I__5277 (
            .O(N__25745),
            .I(N__25727));
    InMux I__5276 (
            .O(N__25744),
            .I(N__25727));
    InMux I__5275 (
            .O(N__25743),
            .I(N__25727));
    InMux I__5274 (
            .O(N__25740),
            .I(N__25722));
    InMux I__5273 (
            .O(N__25739),
            .I(N__25722));
    LocalMux I__5272 (
            .O(N__25736),
            .I(N__25719));
    LocalMux I__5271 (
            .O(N__25727),
            .I(N__25716));
    LocalMux I__5270 (
            .O(N__25722),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.state_1 ));
    Odrv4 I__5269 (
            .O(N__25719),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.state_1 ));
    Odrv4 I__5268 (
            .O(N__25716),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.state_1 ));
    CascadeMux I__5267 (
            .O(N__25709),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n770_cascade_ ));
    InMux I__5266 (
            .O(N__25706),
            .I(N__25703));
    LocalMux I__5265 (
            .O(N__25703),
            .I(N__25700));
    Odrv12 I__5264 (
            .O(N__25700),
            .I(\Inst_core.n6713 ));
    CEMux I__5263 (
            .O(N__25697),
            .I(N__25693));
    CEMux I__5262 (
            .O(N__25696),
            .I(N__25690));
    LocalMux I__5261 (
            .O(N__25693),
            .I(N__25687));
    LocalMux I__5260 (
            .O(N__25690),
            .I(N__25684));
    Span4Mux_v I__5259 (
            .O(N__25687),
            .I(N__25681));
    Span4Mux_h I__5258 (
            .O(N__25684),
            .I(N__25678));
    Odrv4 I__5257 (
            .O(N__25681),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4076 ));
    Odrv4 I__5256 (
            .O(N__25678),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4076 ));
    InMux I__5255 (
            .O(N__25673),
            .I(N__25669));
    InMux I__5254 (
            .O(N__25672),
            .I(N__25666));
    LocalMux I__5253 (
            .O(N__25669),
            .I(N__25663));
    LocalMux I__5252 (
            .O(N__25666),
            .I(configRegister_17_adj_1303));
    Odrv4 I__5251 (
            .O(N__25663),
            .I(configRegister_17_adj_1303));
    InMux I__5250 (
            .O(N__25658),
            .I(N__25655));
    LocalMux I__5249 (
            .O(N__25655),
            .I(N__25652));
    Span4Mux_s2_v I__5248 (
            .O(N__25652),
            .I(N__25648));
    InMux I__5247 (
            .O(N__25651),
            .I(N__25645));
    Odrv4 I__5246 (
            .O(N__25648),
            .I(configRegister_4_adj_1356));
    LocalMux I__5245 (
            .O(N__25645),
            .I(configRegister_4_adj_1356));
    InMux I__5244 (
            .O(N__25640),
            .I(N__25636));
    InMux I__5243 (
            .O(N__25639),
            .I(N__25633));
    LocalMux I__5242 (
            .O(N__25636),
            .I(N__25630));
    LocalMux I__5241 (
            .O(N__25633),
            .I(maskRegister_5_adj_1363));
    Odrv4 I__5240 (
            .O(N__25630),
            .I(maskRegister_5_adj_1363));
    SRMux I__5239 (
            .O(N__25625),
            .I(N__25622));
    LocalMux I__5238 (
            .O(N__25622),
            .I(N__25619));
    Span4Mux_v I__5237 (
            .O(N__25619),
            .I(N__25616));
    Odrv4 I__5236 (
            .O(N__25616),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4764 ));
    CascadeMux I__5235 (
            .O(N__25613),
            .I(N__25610));
    InMux I__5234 (
            .O(N__25610),
            .I(N__25605));
    InMux I__5233 (
            .O(N__25609),
            .I(N__25600));
    InMux I__5232 (
            .O(N__25608),
            .I(N__25600));
    LocalMux I__5231 (
            .O(N__25605),
            .I(N__25594));
    LocalMux I__5230 (
            .O(N__25600),
            .I(N__25594));
    InMux I__5229 (
            .O(N__25599),
            .I(N__25590));
    Span4Mux_v I__5228 (
            .O(N__25594),
            .I(N__25584));
    InMux I__5227 (
            .O(N__25593),
            .I(N__25581));
    LocalMux I__5226 (
            .O(N__25590),
            .I(N__25578));
    InMux I__5225 (
            .O(N__25589),
            .I(N__25571));
    InMux I__5224 (
            .O(N__25588),
            .I(N__25571));
    InMux I__5223 (
            .O(N__25587),
            .I(N__25571));
    Odrv4 I__5222 (
            .O(N__25584),
            .I(cmd_18));
    LocalMux I__5221 (
            .O(N__25581),
            .I(cmd_18));
    Odrv4 I__5220 (
            .O(N__25578),
            .I(cmd_18));
    LocalMux I__5219 (
            .O(N__25571),
            .I(cmd_18));
    InMux I__5218 (
            .O(N__25562),
            .I(N__25559));
    LocalMux I__5217 (
            .O(N__25559),
            .I(N__25555));
    InMux I__5216 (
            .O(N__25558),
            .I(N__25552));
    Odrv4 I__5215 (
            .O(N__25555),
            .I(configRegister_13_adj_1347));
    LocalMux I__5214 (
            .O(N__25552),
            .I(configRegister_13_adj_1347));
    InMux I__5213 (
            .O(N__25547),
            .I(N__25544));
    LocalMux I__5212 (
            .O(N__25544),
            .I(N__25540));
    InMux I__5211 (
            .O(N__25543),
            .I(N__25537));
    Odrv4 I__5210 (
            .O(N__25540),
            .I(configRegister_14_adj_1386));
    LocalMux I__5209 (
            .O(N__25537),
            .I(configRegister_14_adj_1386));
    InMux I__5208 (
            .O(N__25532),
            .I(N__25529));
    LocalMux I__5207 (
            .O(N__25529),
            .I(N__25524));
    InMux I__5206 (
            .O(N__25528),
            .I(N__25519));
    InMux I__5205 (
            .O(N__25527),
            .I(N__25519));
    Odrv4 I__5204 (
            .O(N__25524),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5 ));
    LocalMux I__5203 (
            .O(N__25519),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5 ));
    CascadeMux I__5202 (
            .O(N__25514),
            .I(N__25508));
    InMux I__5201 (
            .O(N__25513),
            .I(N__25504));
    InMux I__5200 (
            .O(N__25512),
            .I(N__25501));
    CascadeMux I__5199 (
            .O(N__25511),
            .I(N__25497));
    InMux I__5198 (
            .O(N__25508),
            .I(N__25494));
    CascadeMux I__5197 (
            .O(N__25507),
            .I(N__25491));
    LocalMux I__5196 (
            .O(N__25504),
            .I(N__25483));
    LocalMux I__5195 (
            .O(N__25501),
            .I(N__25483));
    InMux I__5194 (
            .O(N__25500),
            .I(N__25480));
    InMux I__5193 (
            .O(N__25497),
            .I(N__25477));
    LocalMux I__5192 (
            .O(N__25494),
            .I(N__25474));
    InMux I__5191 (
            .O(N__25491),
            .I(N__25471));
    InMux I__5190 (
            .O(N__25490),
            .I(N__25468));
    InMux I__5189 (
            .O(N__25489),
            .I(N__25465));
    InMux I__5188 (
            .O(N__25488),
            .I(N__25462));
    Span4Mux_v I__5187 (
            .O(N__25483),
            .I(N__25459));
    LocalMux I__5186 (
            .O(N__25480),
            .I(N__25456));
    LocalMux I__5185 (
            .O(N__25477),
            .I(N__25452));
    Span4Mux_v I__5184 (
            .O(N__25474),
            .I(N__25449));
    LocalMux I__5183 (
            .O(N__25471),
            .I(N__25446));
    LocalMux I__5182 (
            .O(N__25468),
            .I(N__25441));
    LocalMux I__5181 (
            .O(N__25465),
            .I(N__25441));
    LocalMux I__5180 (
            .O(N__25462),
            .I(N__25438));
    Span4Mux_v I__5179 (
            .O(N__25459),
            .I(N__25433));
    Span4Mux_v I__5178 (
            .O(N__25456),
            .I(N__25433));
    InMux I__5177 (
            .O(N__25455),
            .I(N__25430));
    Span4Mux_v I__5176 (
            .O(N__25452),
            .I(N__25425));
    Span4Mux_v I__5175 (
            .O(N__25449),
            .I(N__25425));
    Span12Mux_v I__5174 (
            .O(N__25446),
            .I(N__25422));
    Span12Mux_v I__5173 (
            .O(N__25441),
            .I(N__25419));
    Span4Mux_v I__5172 (
            .O(N__25438),
            .I(N__25414));
    Span4Mux_h I__5171 (
            .O(N__25433),
            .I(N__25414));
    LocalMux I__5170 (
            .O(N__25430),
            .I(memoryOut_5));
    Odrv4 I__5169 (
            .O(N__25425),
            .I(memoryOut_5));
    Odrv12 I__5168 (
            .O(N__25422),
            .I(memoryOut_5));
    Odrv12 I__5167 (
            .O(N__25419),
            .I(memoryOut_5));
    Odrv4 I__5166 (
            .O(N__25414),
            .I(memoryOut_5));
    CascadeMux I__5165 (
            .O(N__25403),
            .I(N__25400));
    InMux I__5164 (
            .O(N__25400),
            .I(N__25394));
    InMux I__5163 (
            .O(N__25399),
            .I(N__25394));
    LocalMux I__5162 (
            .O(N__25394),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n554 ));
    CascadeMux I__5161 (
            .O(N__25391),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n22_cascade_ ));
    CascadeMux I__5160 (
            .O(N__25388),
            .I(\Inst_core.n8515_cascade_ ));
    InMux I__5159 (
            .O(N__25385),
            .I(N__25379));
    InMux I__5158 (
            .O(N__25384),
            .I(N__25379));
    LocalMux I__5157 (
            .O(N__25379),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n451 ));
    InMux I__5156 (
            .O(N__25376),
            .I(N__25370));
    InMux I__5155 (
            .O(N__25375),
            .I(N__25370));
    LocalMux I__5154 (
            .O(N__25370),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n760 ));
    InMux I__5153 (
            .O(N__25367),
            .I(N__25358));
    InMux I__5152 (
            .O(N__25366),
            .I(N__25349));
    InMux I__5151 (
            .O(N__25365),
            .I(N__25349));
    InMux I__5150 (
            .O(N__25364),
            .I(N__25349));
    InMux I__5149 (
            .O(N__25363),
            .I(N__25349));
    InMux I__5148 (
            .O(N__25362),
            .I(N__25344));
    InMux I__5147 (
            .O(N__25361),
            .I(N__25344));
    LocalMux I__5146 (
            .O(N__25358),
            .I(N__25341));
    LocalMux I__5145 (
            .O(N__25349),
            .I(N__25338));
    LocalMux I__5144 (
            .O(N__25344),
            .I(N__25331));
    Span4Mux_v I__5143 (
            .O(N__25341),
            .I(N__25331));
    Span4Mux_s2_v I__5142 (
            .O(N__25338),
            .I(N__25331));
    Odrv4 I__5141 (
            .O(N__25331),
            .I(\Inst_core.n31 ));
    CascadeMux I__5140 (
            .O(N__25328),
            .I(N__25317));
    CascadeMux I__5139 (
            .O(N__25327),
            .I(N__25313));
    CascadeMux I__5138 (
            .O(N__25326),
            .I(N__25309));
    CascadeMux I__5137 (
            .O(N__25325),
            .I(N__25305));
    CascadeMux I__5136 (
            .O(N__25324),
            .I(N__25302));
    CascadeMux I__5135 (
            .O(N__25323),
            .I(N__25298));
    CascadeMux I__5134 (
            .O(N__25322),
            .I(N__25294));
    CascadeMux I__5133 (
            .O(N__25321),
            .I(N__25290));
    InMux I__5132 (
            .O(N__25320),
            .I(N__25273));
    InMux I__5131 (
            .O(N__25317),
            .I(N__25273));
    InMux I__5130 (
            .O(N__25316),
            .I(N__25273));
    InMux I__5129 (
            .O(N__25313),
            .I(N__25273));
    InMux I__5128 (
            .O(N__25312),
            .I(N__25273));
    InMux I__5127 (
            .O(N__25309),
            .I(N__25273));
    InMux I__5126 (
            .O(N__25308),
            .I(N__25273));
    InMux I__5125 (
            .O(N__25305),
            .I(N__25273));
    InMux I__5124 (
            .O(N__25302),
            .I(N__25258));
    InMux I__5123 (
            .O(N__25301),
            .I(N__25258));
    InMux I__5122 (
            .O(N__25298),
            .I(N__25258));
    InMux I__5121 (
            .O(N__25297),
            .I(N__25258));
    InMux I__5120 (
            .O(N__25294),
            .I(N__25258));
    InMux I__5119 (
            .O(N__25293),
            .I(N__25258));
    InMux I__5118 (
            .O(N__25290),
            .I(N__25258));
    LocalMux I__5117 (
            .O(N__25273),
            .I(N__25255));
    LocalMux I__5116 (
            .O(N__25258),
            .I(N__25252));
    Span4Mux_h I__5115 (
            .O(N__25255),
            .I(N__25249));
    Span4Mux_h I__5114 (
            .O(N__25252),
            .I(N__25246));
    Odrv4 I__5113 (
            .O(N__25249),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n1765 ));
    Odrv4 I__5112 (
            .O(N__25246),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n1765 ));
    InMux I__5111 (
            .O(N__25241),
            .I(N__25238));
    LocalMux I__5110 (
            .O(N__25238),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n667 ));
    CascadeMux I__5109 (
            .O(N__25235),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n667_cascade_ ));
    InMux I__5108 (
            .O(N__25232),
            .I(N__25229));
    LocalMux I__5107 (
            .O(N__25229),
            .I(N__25222));
    InMux I__5106 (
            .O(N__25228),
            .I(N__25213));
    InMux I__5105 (
            .O(N__25227),
            .I(N__25213));
    InMux I__5104 (
            .O(N__25226),
            .I(N__25213));
    InMux I__5103 (
            .O(N__25225),
            .I(N__25213));
    Odrv4 I__5102 (
            .O(N__25222),
            .I(\Inst_core.n31_adj_1174 ));
    LocalMux I__5101 (
            .O(N__25213),
            .I(\Inst_core.n31_adj_1174 ));
    CascadeMux I__5100 (
            .O(N__25208),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n100_cascade_ ));
    InMux I__5099 (
            .O(N__25205),
            .I(N__25199));
    InMux I__5098 (
            .O(N__25204),
            .I(N__25199));
    LocalMux I__5097 (
            .O(N__25199),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n656 ));
    InMux I__5096 (
            .O(N__25196),
            .I(N__25193));
    LocalMux I__5095 (
            .O(N__25193),
            .I(\Inst_core.n8518 ));
    CascadeMux I__5094 (
            .O(N__25190),
            .I(N__25187));
    InMux I__5093 (
            .O(N__25187),
            .I(N__25179));
    InMux I__5092 (
            .O(N__25186),
            .I(N__25176));
    InMux I__5091 (
            .O(N__25185),
            .I(N__25173));
    InMux I__5090 (
            .O(N__25184),
            .I(N__25170));
    InMux I__5089 (
            .O(N__25183),
            .I(N__25165));
    InMux I__5088 (
            .O(N__25182),
            .I(N__25165));
    LocalMux I__5087 (
            .O(N__25179),
            .I(\Inst_core.state_1_adj_1134 ));
    LocalMux I__5086 (
            .O(N__25176),
            .I(\Inst_core.state_1_adj_1134 ));
    LocalMux I__5085 (
            .O(N__25173),
            .I(\Inst_core.state_1_adj_1134 ));
    LocalMux I__5084 (
            .O(N__25170),
            .I(\Inst_core.state_1_adj_1134 ));
    LocalMux I__5083 (
            .O(N__25165),
            .I(\Inst_core.state_1_adj_1134 ));
    InMux I__5082 (
            .O(N__25154),
            .I(N__25148));
    InMux I__5081 (
            .O(N__25153),
            .I(N__25148));
    LocalMux I__5080 (
            .O(N__25148),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n657 ));
    InMux I__5079 (
            .O(N__25145),
            .I(N__25141));
    CascadeMux I__5078 (
            .O(N__25144),
            .I(N__25138));
    LocalMux I__5077 (
            .O(N__25141),
            .I(N__25134));
    InMux I__5076 (
            .O(N__25138),
            .I(N__25129));
    InMux I__5075 (
            .O(N__25137),
            .I(N__25129));
    Odrv4 I__5074 (
            .O(N__25134),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4 ));
    LocalMux I__5073 (
            .O(N__25129),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4 ));
    InMux I__5072 (
            .O(N__25124),
            .I(N__25121));
    LocalMux I__5071 (
            .O(N__25121),
            .I(N__25116));
    InMux I__5070 (
            .O(N__25120),
            .I(N__25111));
    InMux I__5069 (
            .O(N__25119),
            .I(N__25111));
    Odrv4 I__5068 (
            .O(N__25116),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5 ));
    LocalMux I__5067 (
            .O(N__25111),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5 ));
    CascadeMux I__5066 (
            .O(N__25106),
            .I(N__25103));
    InMux I__5065 (
            .O(N__25103),
            .I(N__25100));
    LocalMux I__5064 (
            .O(N__25100),
            .I(N__25097));
    Span4Mux_v I__5063 (
            .O(N__25097),
            .I(N__25094));
    Odrv4 I__5062 (
            .O(N__25094),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_7 ));
    CascadeMux I__5061 (
            .O(N__25091),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n8844_cascade_ ));
    InMux I__5060 (
            .O(N__25088),
            .I(N__25085));
    LocalMux I__5059 (
            .O(N__25085),
            .I(\Inst_core.Inst_decoder.n6 ));
    InMux I__5058 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__5057 (
            .O(N__25079),
            .I(N__25076));
    Span4Mux_h I__5056 (
            .O(N__25076),
            .I(N__25073));
    Odrv4 I__5055 (
            .O(N__25073),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9052 ));
    InMux I__5054 (
            .O(N__25070),
            .I(N__25067));
    LocalMux I__5053 (
            .O(N__25067),
            .I(N__25063));
    InMux I__5052 (
            .O(N__25066),
            .I(N__25060));
    Odrv12 I__5051 (
            .O(N__25063),
            .I(valueRegister_1_adj_1335));
    LocalMux I__5050 (
            .O(N__25060),
            .I(valueRegister_1_adj_1335));
    InMux I__5049 (
            .O(N__25055),
            .I(N__25051));
    InMux I__5048 (
            .O(N__25054),
            .I(N__25047));
    LocalMux I__5047 (
            .O(N__25051),
            .I(N__25044));
    InMux I__5046 (
            .O(N__25050),
            .I(N__25041));
    LocalMux I__5045 (
            .O(N__25047),
            .I(N__25036));
    Span4Mux_s3_v I__5044 (
            .O(N__25044),
            .I(N__25036));
    LocalMux I__5043 (
            .O(N__25041),
            .I(divider_20));
    Odrv4 I__5042 (
            .O(N__25036),
            .I(divider_20));
    CascadeMux I__5041 (
            .O(N__25031),
            .I(N__25028));
    InMux I__5040 (
            .O(N__25028),
            .I(N__25024));
    InMux I__5039 (
            .O(N__25027),
            .I(N__25020));
    LocalMux I__5038 (
            .O(N__25024),
            .I(N__25017));
    InMux I__5037 (
            .O(N__25023),
            .I(N__25014));
    LocalMux I__5036 (
            .O(N__25020),
            .I(divider_21));
    Odrv4 I__5035 (
            .O(N__25017),
            .I(divider_21));
    LocalMux I__5034 (
            .O(N__25014),
            .I(divider_21));
    InMux I__5033 (
            .O(N__25007),
            .I(N__25004));
    LocalMux I__5032 (
            .O(N__25004),
            .I(N__25001));
    Odrv4 I__5031 (
            .O(N__25001),
            .I(\Inst_core.Inst_sampler.n8598 ));
    InMux I__5030 (
            .O(N__24998),
            .I(N__24995));
    LocalMux I__5029 (
            .O(N__24995),
            .I(N__24992));
    Odrv4 I__5028 (
            .O(N__24992),
            .I(\Inst_core.Inst_sampler.n8602 ));
    CascadeMux I__5027 (
            .O(N__24989),
            .I(\Inst_core.Inst_sampler.n8600_cascade_ ));
    InMux I__5026 (
            .O(N__24986),
            .I(N__24983));
    LocalMux I__5025 (
            .O(N__24983),
            .I(\Inst_core.Inst_sampler.n8604 ));
    CascadeMux I__5024 (
            .O(N__24980),
            .I(N__24977));
    InMux I__5023 (
            .O(N__24977),
            .I(N__24974));
    LocalMux I__5022 (
            .O(N__24974),
            .I(N__24970));
    InMux I__5021 (
            .O(N__24973),
            .I(N__24967));
    Span4Mux_s3_v I__5020 (
            .O(N__24970),
            .I(N__24964));
    LocalMux I__5019 (
            .O(N__24967),
            .I(N__24959));
    Span4Mux_v I__5018 (
            .O(N__24964),
            .I(N__24959));
    Odrv4 I__5017 (
            .O(N__24959),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelL16 ));
    InMux I__5016 (
            .O(N__24956),
            .I(N__24953));
    LocalMux I__5015 (
            .O(N__24953),
            .I(N__24950));
    Span12Mux_s6_h I__5014 (
            .O(N__24950),
            .I(N__24946));
    InMux I__5013 (
            .O(N__24949),
            .I(N__24943));
    Odrv12 I__5012 (
            .O(N__24946),
            .I(configRegister_24_adj_1338));
    LocalMux I__5011 (
            .O(N__24943),
            .I(configRegister_24_adj_1338));
    InMux I__5010 (
            .O(N__24938),
            .I(N__24932));
    InMux I__5009 (
            .O(N__24937),
            .I(N__24932));
    LocalMux I__5008 (
            .O(N__24932),
            .I(N__24929));
    Span4Mux_h I__5007 (
            .O(N__24929),
            .I(N__24925));
    InMux I__5006 (
            .O(N__24928),
            .I(N__24922));
    Span4Mux_v I__5005 (
            .O(N__24925),
            .I(N__24919));
    LocalMux I__5004 (
            .O(N__24922),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16 ));
    Odrv4 I__5003 (
            .O(N__24919),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16 ));
    InMux I__5002 (
            .O(N__24914),
            .I(N__24909));
    InMux I__5001 (
            .O(N__24913),
            .I(N__24904));
    InMux I__5000 (
            .O(N__24912),
            .I(N__24904));
    LocalMux I__4999 (
            .O(N__24909),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1 ));
    LocalMux I__4998 (
            .O(N__24904),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1 ));
    CascadeMux I__4997 (
            .O(N__24899),
            .I(N__24896));
    InMux I__4996 (
            .O(N__24896),
            .I(N__24892));
    InMux I__4995 (
            .O(N__24895),
            .I(N__24889));
    LocalMux I__4994 (
            .O(N__24892),
            .I(N__24883));
    LocalMux I__4993 (
            .O(N__24889),
            .I(N__24883));
    InMux I__4992 (
            .O(N__24888),
            .I(N__24880));
    Span4Mux_v I__4991 (
            .O(N__24883),
            .I(N__24877));
    LocalMux I__4990 (
            .O(N__24880),
            .I(divider_9));
    Odrv4 I__4989 (
            .O(N__24877),
            .I(divider_9));
    CascadeMux I__4988 (
            .O(N__24872),
            .I(N__24868));
    InMux I__4987 (
            .O(N__24871),
            .I(N__24864));
    InMux I__4986 (
            .O(N__24868),
            .I(N__24861));
    InMux I__4985 (
            .O(N__24867),
            .I(N__24858));
    LocalMux I__4984 (
            .O(N__24864),
            .I(N__24853));
    LocalMux I__4983 (
            .O(N__24861),
            .I(N__24853));
    LocalMux I__4982 (
            .O(N__24858),
            .I(divider_7));
    Odrv4 I__4981 (
            .O(N__24853),
            .I(divider_7));
    InMux I__4980 (
            .O(N__24848),
            .I(N__24845));
    LocalMux I__4979 (
            .O(N__24845),
            .I(\Inst_core.Inst_sampler.n29 ));
    InMux I__4978 (
            .O(N__24842),
            .I(N__24839));
    LocalMux I__4977 (
            .O(N__24839),
            .I(N__24836));
    Odrv4 I__4976 (
            .O(N__24836),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_7 ));
    InMux I__4975 (
            .O(N__24833),
            .I(N__24830));
    LocalMux I__4974 (
            .O(N__24830),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_4 ));
    InMux I__4973 (
            .O(N__24827),
            .I(N__24824));
    LocalMux I__4972 (
            .O(N__24824),
            .I(N__24820));
    InMux I__4971 (
            .O(N__24823),
            .I(N__24817));
    Odrv4 I__4970 (
            .O(N__24820),
            .I(valueRegister_5_adj_1331));
    LocalMux I__4969 (
            .O(N__24817),
            .I(valueRegister_5_adj_1331));
    CascadeMux I__4968 (
            .O(N__24812),
            .I(N__24809));
    InMux I__4967 (
            .O(N__24809),
            .I(N__24806));
    LocalMux I__4966 (
            .O(N__24806),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_5 ));
    InMux I__4965 (
            .O(N__24803),
            .I(N__24798));
    InMux I__4964 (
            .O(N__24802),
            .I(N__24795));
    InMux I__4963 (
            .O(N__24801),
            .I(N__24792));
    LocalMux I__4962 (
            .O(N__24798),
            .I(divider_15));
    LocalMux I__4961 (
            .O(N__24795),
            .I(divider_15));
    LocalMux I__4960 (
            .O(N__24792),
            .I(divider_15));
    CascadeMux I__4959 (
            .O(N__24785),
            .I(N__24782));
    InMux I__4958 (
            .O(N__24782),
            .I(N__24779));
    LocalMux I__4957 (
            .O(N__24779),
            .I(N__24775));
    CascadeMux I__4956 (
            .O(N__24778),
            .I(N__24772));
    Span4Mux_h I__4955 (
            .O(N__24775),
            .I(N__24768));
    InMux I__4954 (
            .O(N__24772),
            .I(N__24765));
    InMux I__4953 (
            .O(N__24771),
            .I(N__24762));
    Span4Mux_v I__4952 (
            .O(N__24768),
            .I(N__24759));
    LocalMux I__4951 (
            .O(N__24765),
            .I(N__24756));
    LocalMux I__4950 (
            .O(N__24762),
            .I(divider_13));
    Odrv4 I__4949 (
            .O(N__24759),
            .I(divider_13));
    Odrv12 I__4948 (
            .O(N__24756),
            .I(divider_13));
    InMux I__4947 (
            .O(N__24749),
            .I(N__24744));
    InMux I__4946 (
            .O(N__24748),
            .I(N__24741));
    InMux I__4945 (
            .O(N__24747),
            .I(N__24738));
    LocalMux I__4944 (
            .O(N__24744),
            .I(divider_16));
    LocalMux I__4943 (
            .O(N__24741),
            .I(divider_16));
    LocalMux I__4942 (
            .O(N__24738),
            .I(divider_16));
    InMux I__4941 (
            .O(N__24731),
            .I(N__24728));
    LocalMux I__4940 (
            .O(N__24728),
            .I(\Inst_core.Inst_sampler.n32 ));
    CascadeMux I__4939 (
            .O(N__24725),
            .I(N__24721));
    CascadeMux I__4938 (
            .O(N__24724),
            .I(N__24718));
    InMux I__4937 (
            .O(N__24721),
            .I(N__24715));
    InMux I__4936 (
            .O(N__24718),
            .I(N__24712));
    LocalMux I__4935 (
            .O(N__24715),
            .I(N__24706));
    LocalMux I__4934 (
            .O(N__24712),
            .I(N__24706));
    InMux I__4933 (
            .O(N__24711),
            .I(N__24703));
    Span4Mux_v I__4932 (
            .O(N__24706),
            .I(N__24700));
    LocalMux I__4931 (
            .O(N__24703),
            .I(divider_14));
    Odrv4 I__4930 (
            .O(N__24700),
            .I(divider_14));
    CascadeMux I__4929 (
            .O(N__24695),
            .I(\Inst_core.Inst_sampler.n8596_cascade_ ));
    InMux I__4928 (
            .O(N__24692),
            .I(N__24689));
    LocalMux I__4927 (
            .O(N__24689),
            .I(\Inst_core.Inst_sampler.n8590 ));
    InMux I__4926 (
            .O(N__24686),
            .I(N__24681));
    InMux I__4925 (
            .O(N__24685),
            .I(N__24678));
    CascadeMux I__4924 (
            .O(N__24684),
            .I(N__24675));
    LocalMux I__4923 (
            .O(N__24681),
            .I(N__24670));
    LocalMux I__4922 (
            .O(N__24678),
            .I(N__24670));
    InMux I__4921 (
            .O(N__24675),
            .I(N__24665));
    Span4Mux_v I__4920 (
            .O(N__24670),
            .I(N__24659));
    InMux I__4919 (
            .O(N__24669),
            .I(N__24654));
    InMux I__4918 (
            .O(N__24668),
            .I(N__24654));
    LocalMux I__4917 (
            .O(N__24665),
            .I(N__24651));
    InMux I__4916 (
            .O(N__24664),
            .I(N__24644));
    InMux I__4915 (
            .O(N__24663),
            .I(N__24644));
    InMux I__4914 (
            .O(N__24662),
            .I(N__24644));
    Odrv4 I__4913 (
            .O(N__24659),
            .I(cmd_29));
    LocalMux I__4912 (
            .O(N__24654),
            .I(cmd_29));
    Odrv4 I__4911 (
            .O(N__24651),
            .I(cmd_29));
    LocalMux I__4910 (
            .O(N__24644),
            .I(cmd_29));
    InMux I__4909 (
            .O(N__24635),
            .I(N__24632));
    LocalMux I__4908 (
            .O(N__24632),
            .I(syncedInput_0));
    CascadeMux I__4907 (
            .O(N__24629),
            .I(N__24626));
    InMux I__4906 (
            .O(N__24626),
            .I(N__24623));
    LocalMux I__4905 (
            .O(N__24623),
            .I(N__24620));
    Span4Mux_v I__4904 (
            .O(N__24620),
            .I(N__24617));
    Odrv4 I__4903 (
            .O(N__24617),
            .I(syncedInput_1));
    CascadeMux I__4902 (
            .O(N__24614),
            .I(N__24611));
    InMux I__4901 (
            .O(N__24611),
            .I(N__24608));
    LocalMux I__4900 (
            .O(N__24608),
            .I(N__24604));
    InMux I__4899 (
            .O(N__24607),
            .I(N__24601));
    Odrv4 I__4898 (
            .O(N__24604),
            .I(valueRegister_4_adj_1332));
    LocalMux I__4897 (
            .O(N__24601),
            .I(valueRegister_4_adj_1332));
    SRMux I__4896 (
            .O(N__24596),
            .I(N__24593));
    LocalMux I__4895 (
            .O(N__24593),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4756 ));
    CascadeMux I__4894 (
            .O(N__24590),
            .I(\Inst_core.Inst_sampler.n31_adj_995_cascade_ ));
    InMux I__4893 (
            .O(N__24587),
            .I(N__24584));
    LocalMux I__4892 (
            .O(N__24584),
            .I(N__24581));
    Span4Mux_h I__4891 (
            .O(N__24581),
            .I(N__24577));
    CascadeMux I__4890 (
            .O(N__24580),
            .I(N__24574));
    Span4Mux_v I__4889 (
            .O(N__24577),
            .I(N__24570));
    InMux I__4888 (
            .O(N__24574),
            .I(N__24565));
    InMux I__4887 (
            .O(N__24573),
            .I(N__24565));
    Odrv4 I__4886 (
            .O(N__24570),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4 ));
    LocalMux I__4885 (
            .O(N__24565),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4 ));
    CascadeMux I__4884 (
            .O(N__24560),
            .I(N__24557));
    InMux I__4883 (
            .O(N__24557),
            .I(N__24554));
    LocalMux I__4882 (
            .O(N__24554),
            .I(N__24551));
    Span4Mux_h I__4881 (
            .O(N__24551),
            .I(N__24547));
    InMux I__4880 (
            .O(N__24550),
            .I(N__24544));
    Odrv4 I__4879 (
            .O(N__24547),
            .I(valueRegister_4_adj_1292));
    LocalMux I__4878 (
            .O(N__24544),
            .I(valueRegister_4_adj_1292));
    SRMux I__4877 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__4876 (
            .O(N__24536),
            .I(N__24533));
    Span4Mux_v I__4875 (
            .O(N__24533),
            .I(N__24530));
    Odrv4 I__4874 (
            .O(N__24530),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4749 ));
    InMux I__4873 (
            .O(N__24527),
            .I(N__24524));
    LocalMux I__4872 (
            .O(N__24524),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_5 ));
    CascadeMux I__4871 (
            .O(N__24521),
            .I(N__24518));
    InMux I__4870 (
            .O(N__24518),
            .I(N__24515));
    LocalMux I__4869 (
            .O(N__24515),
            .I(N__24512));
    Odrv12 I__4868 (
            .O(N__24512),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_7 ));
    InMux I__4867 (
            .O(N__24509),
            .I(N__24506));
    LocalMux I__4866 (
            .O(N__24506),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_4 ));
    InMux I__4865 (
            .O(N__24503),
            .I(N__24499));
    InMux I__4864 (
            .O(N__24502),
            .I(N__24496));
    LocalMux I__4863 (
            .O(N__24499),
            .I(N__24493));
    LocalMux I__4862 (
            .O(N__24496),
            .I(fwd_12));
    Odrv4 I__4861 (
            .O(N__24493),
            .I(fwd_12));
    CascadeMux I__4860 (
            .O(N__24488),
            .I(N__24485));
    InMux I__4859 (
            .O(N__24485),
            .I(N__24481));
    InMux I__4858 (
            .O(N__24484),
            .I(N__24478));
    LocalMux I__4857 (
            .O(N__24481),
            .I(N__24475));
    LocalMux I__4856 (
            .O(N__24478),
            .I(fwd_1));
    Odrv4 I__4855 (
            .O(N__24475),
            .I(fwd_1));
    InMux I__4854 (
            .O(N__24470),
            .I(N__24467));
    LocalMux I__4853 (
            .O(N__24467),
            .I(\Inst_core.Inst_controller.n13 ));
    InMux I__4852 (
            .O(N__24464),
            .I(N__24460));
    InMux I__4851 (
            .O(N__24463),
            .I(N__24457));
    LocalMux I__4850 (
            .O(N__24460),
            .I(N__24454));
    LocalMux I__4849 (
            .O(N__24457),
            .I(bwd_10));
    Odrv12 I__4848 (
            .O(N__24454),
            .I(bwd_10));
    InMux I__4847 (
            .O(N__24449),
            .I(N__24446));
    LocalMux I__4846 (
            .O(N__24446),
            .I(\Inst_core.Inst_controller.n14 ));
    InMux I__4845 (
            .O(N__24443),
            .I(N__24440));
    LocalMux I__4844 (
            .O(N__24440),
            .I(N__24437));
    Span4Mux_v I__4843 (
            .O(N__24437),
            .I(N__24433));
    InMux I__4842 (
            .O(N__24436),
            .I(N__24430));
    Sp12to4 I__4841 (
            .O(N__24433),
            .I(N__24427));
    LocalMux I__4840 (
            .O(N__24430),
            .I(fwd_8));
    Odrv12 I__4839 (
            .O(N__24427),
            .I(fwd_8));
    InMux I__4838 (
            .O(N__24422),
            .I(N__24419));
    LocalMux I__4837 (
            .O(N__24419),
            .I(\Inst_core.Inst_controller.n11 ));
    InMux I__4836 (
            .O(N__24416),
            .I(N__24413));
    LocalMux I__4835 (
            .O(N__24413),
            .I(N__24410));
    Span4Mux_h I__4834 (
            .O(N__24410),
            .I(N__24407));
    Span4Mux_h I__4833 (
            .O(N__24407),
            .I(N__24404));
    Odrv4 I__4832 (
            .O(N__24404),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n14 ));
    InMux I__4831 (
            .O(N__24401),
            .I(N__24398));
    LocalMux I__4830 (
            .O(N__24398),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n11 ));
    CascadeMux I__4829 (
            .O(N__24395),
            .I(N__24392));
    InMux I__4828 (
            .O(N__24392),
            .I(N__24385));
    InMux I__4827 (
            .O(N__24391),
            .I(N__24385));
    CascadeMux I__4826 (
            .O(N__24390),
            .I(N__24382));
    LocalMux I__4825 (
            .O(N__24385),
            .I(N__24379));
    InMux I__4824 (
            .O(N__24382),
            .I(N__24376));
    Odrv4 I__4823 (
            .O(N__24379),
            .I(cmd_37));
    LocalMux I__4822 (
            .O(N__24376),
            .I(cmd_37));
    InMux I__4821 (
            .O(N__24371),
            .I(N__24368));
    LocalMux I__4820 (
            .O(N__24368),
            .I(N__24363));
    InMux I__4819 (
            .O(N__24367),
            .I(N__24358));
    InMux I__4818 (
            .O(N__24366),
            .I(N__24358));
    Odrv4 I__4817 (
            .O(N__24363),
            .I(cmd_36));
    LocalMux I__4816 (
            .O(N__24358),
            .I(cmd_36));
    InMux I__4815 (
            .O(N__24353),
            .I(N__24350));
    LocalMux I__4814 (
            .O(N__24350),
            .I(N__24347));
    Span12Mux_s3_v I__4813 (
            .O(N__24347),
            .I(N__24343));
    InMux I__4812 (
            .O(N__24346),
            .I(N__24340));
    Odrv12 I__4811 (
            .O(N__24343),
            .I(configRegister_6_adj_1354));
    LocalMux I__4810 (
            .O(N__24340),
            .I(configRegister_6_adj_1354));
    InMux I__4809 (
            .O(N__24335),
            .I(N__24332));
    LocalMux I__4808 (
            .O(N__24332),
            .I(N__24329));
    Span4Mux_h I__4807 (
            .O(N__24329),
            .I(N__24325));
    InMux I__4806 (
            .O(N__24328),
            .I(N__24322));
    Odrv4 I__4805 (
            .O(N__24325),
            .I(valueRegister_5_adj_1291));
    LocalMux I__4804 (
            .O(N__24322),
            .I(valueRegister_5_adj_1291));
    InMux I__4803 (
            .O(N__24317),
            .I(N__24314));
    LocalMux I__4802 (
            .O(N__24314),
            .I(N__24311));
    Span4Mux_h I__4801 (
            .O(N__24311),
            .I(N__24306));
    InMux I__4800 (
            .O(N__24310),
            .I(N__24301));
    InMux I__4799 (
            .O(N__24309),
            .I(N__24301));
    Odrv4 I__4798 (
            .O(N__24306),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5 ));
    LocalMux I__4797 (
            .O(N__24301),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5 ));
    SRMux I__4796 (
            .O(N__24296),
            .I(N__24293));
    LocalMux I__4795 (
            .O(N__24293),
            .I(N__24290));
    Span4Mux_h I__4794 (
            .O(N__24290),
            .I(N__24287));
    Odrv4 I__4793 (
            .O(N__24287),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4750 ));
    InMux I__4792 (
            .O(N__24284),
            .I(N__24280));
    InMux I__4791 (
            .O(N__24283),
            .I(N__24277));
    LocalMux I__4790 (
            .O(N__24280),
            .I(N__24274));
    LocalMux I__4789 (
            .O(N__24277),
            .I(bwd_11));
    Odrv12 I__4788 (
            .O(N__24274),
            .I(bwd_11));
    CascadeMux I__4787 (
            .O(N__24269),
            .I(N__24266));
    InMux I__4786 (
            .O(N__24266),
            .I(N__24262));
    InMux I__4785 (
            .O(N__24265),
            .I(N__24259));
    LocalMux I__4784 (
            .O(N__24262),
            .I(N__24256));
    LocalMux I__4783 (
            .O(N__24259),
            .I(bwd_8));
    Odrv4 I__4782 (
            .O(N__24256),
            .I(bwd_8));
    InMux I__4781 (
            .O(N__24251),
            .I(N__24247));
    InMux I__4780 (
            .O(N__24250),
            .I(N__24244));
    LocalMux I__4779 (
            .O(N__24247),
            .I(fwd_11));
    LocalMux I__4778 (
            .O(N__24244),
            .I(fwd_11));
    CascadeMux I__4777 (
            .O(N__24239),
            .I(N__24236));
    InMux I__4776 (
            .O(N__24236),
            .I(N__24232));
    InMux I__4775 (
            .O(N__24235),
            .I(N__24229));
    LocalMux I__4774 (
            .O(N__24232),
            .I(N__24224));
    LocalMux I__4773 (
            .O(N__24229),
            .I(N__24224));
    Odrv4 I__4772 (
            .O(N__24224),
            .I(fwd_4));
    CascadeMux I__4771 (
            .O(N__24221),
            .I(\Inst_core.Inst_controller.n18_cascade_ ));
    InMux I__4770 (
            .O(N__24218),
            .I(N__24215));
    LocalMux I__4769 (
            .O(N__24215),
            .I(\Inst_core.Inst_controller.n21 ));
    InMux I__4768 (
            .O(N__24212),
            .I(N__24208));
    InMux I__4767 (
            .O(N__24211),
            .I(N__24205));
    LocalMux I__4766 (
            .O(N__24208),
            .I(fwd_13));
    LocalMux I__4765 (
            .O(N__24205),
            .I(fwd_13));
    CascadeMux I__4764 (
            .O(N__24200),
            .I(N__24196));
    InMux I__4763 (
            .O(N__24199),
            .I(N__24193));
    InMux I__4762 (
            .O(N__24196),
            .I(N__24190));
    LocalMux I__4761 (
            .O(N__24193),
            .I(fwd_9));
    LocalMux I__4760 (
            .O(N__24190),
            .I(fwd_9));
    InMux I__4759 (
            .O(N__24185),
            .I(N__24182));
    LocalMux I__4758 (
            .O(N__24182),
            .I(\Inst_core.Inst_controller.n15 ));
    InMux I__4757 (
            .O(N__24179),
            .I(N__24172));
    CascadeMux I__4756 (
            .O(N__24178),
            .I(N__24169));
    InMux I__4755 (
            .O(N__24177),
            .I(N__24163));
    InMux I__4754 (
            .O(N__24176),
            .I(N__24163));
    InMux I__4753 (
            .O(N__24175),
            .I(N__24160));
    LocalMux I__4752 (
            .O(N__24172),
            .I(N__24157));
    InMux I__4751 (
            .O(N__24169),
            .I(N__24154));
    CascadeMux I__4750 (
            .O(N__24168),
            .I(N__24149));
    LocalMux I__4749 (
            .O(N__24163),
            .I(N__24146));
    LocalMux I__4748 (
            .O(N__24160),
            .I(N__24143));
    Span4Mux_v I__4747 (
            .O(N__24157),
            .I(N__24138));
    LocalMux I__4746 (
            .O(N__24154),
            .I(N__24138));
    InMux I__4745 (
            .O(N__24153),
            .I(N__24135));
    InMux I__4744 (
            .O(N__24152),
            .I(N__24130));
    InMux I__4743 (
            .O(N__24149),
            .I(N__24130));
    Odrv4 I__4742 (
            .O(N__24146),
            .I(cmd_30));
    Odrv4 I__4741 (
            .O(N__24143),
            .I(cmd_30));
    Odrv4 I__4740 (
            .O(N__24138),
            .I(cmd_30));
    LocalMux I__4739 (
            .O(N__24135),
            .I(cmd_30));
    LocalMux I__4738 (
            .O(N__24130),
            .I(cmd_30));
    InMux I__4737 (
            .O(N__24119),
            .I(N__24112));
    InMux I__4736 (
            .O(N__24118),
            .I(N__24112));
    InMux I__4735 (
            .O(N__24117),
            .I(N__24109));
    LocalMux I__4734 (
            .O(N__24112),
            .I(N__24106));
    LocalMux I__4733 (
            .O(N__24109),
            .I(configRegister_22));
    Odrv12 I__4732 (
            .O(N__24106),
            .I(configRegister_22));
    InMux I__4731 (
            .O(N__24101),
            .I(N__24096));
    InMux I__4730 (
            .O(N__24100),
            .I(N__24093));
    InMux I__4729 (
            .O(N__24099),
            .I(N__24090));
    LocalMux I__4728 (
            .O(N__24096),
            .I(cmd_33));
    LocalMux I__4727 (
            .O(N__24093),
            .I(cmd_33));
    LocalMux I__4726 (
            .O(N__24090),
            .I(cmd_33));
    InMux I__4725 (
            .O(N__24083),
            .I(N__24080));
    LocalMux I__4724 (
            .O(N__24080),
            .I(N__24077));
    Span4Mux_v I__4723 (
            .O(N__24077),
            .I(N__24074));
    Span4Mux_h I__4722 (
            .O(N__24074),
            .I(N__24070));
    InMux I__4721 (
            .O(N__24073),
            .I(N__24067));
    Odrv4 I__4720 (
            .O(N__24070),
            .I(configRegister_9_adj_1391));
    LocalMux I__4719 (
            .O(N__24067),
            .I(configRegister_9_adj_1391));
    InMux I__4718 (
            .O(N__24062),
            .I(N__24058));
    InMux I__4717 (
            .O(N__24061),
            .I(N__24055));
    LocalMux I__4716 (
            .O(N__24058),
            .I(N__24050));
    LocalMux I__4715 (
            .O(N__24055),
            .I(N__24050));
    Span4Mux_v I__4714 (
            .O(N__24050),
            .I(N__24046));
    InMux I__4713 (
            .O(N__24049),
            .I(N__24043));
    Span4Mux_h I__4712 (
            .O(N__24046),
            .I(N__24040));
    LocalMux I__4711 (
            .O(N__24043),
            .I(cmd_38));
    Odrv4 I__4710 (
            .O(N__24040),
            .I(cmd_38));
    InMux I__4709 (
            .O(N__24035),
            .I(N__24031));
    InMux I__4708 (
            .O(N__24034),
            .I(N__24028));
    LocalMux I__4707 (
            .O(N__24031),
            .I(N__24025));
    LocalMux I__4706 (
            .O(N__24028),
            .I(N__24020));
    Span4Mux_v I__4705 (
            .O(N__24025),
            .I(N__24020));
    Odrv4 I__4704 (
            .O(N__24020),
            .I(\Inst_core.Inst_controller.fwd_14 ));
    InMux I__4703 (
            .O(N__24017),
            .I(N__24014));
    LocalMux I__4702 (
            .O(N__24014),
            .I(N__24011));
    Span4Mux_s2_v I__4701 (
            .O(N__24011),
            .I(N__24007));
    InMux I__4700 (
            .O(N__24010),
            .I(N__24004));
    Odrv4 I__4699 (
            .O(N__24007),
            .I(configRegister_8_adj_1352));
    LocalMux I__4698 (
            .O(N__24004),
            .I(configRegister_8_adj_1352));
    InMux I__4697 (
            .O(N__23999),
            .I(N__23994));
    InMux I__4696 (
            .O(N__23998),
            .I(N__23989));
    InMux I__4695 (
            .O(N__23997),
            .I(N__23986));
    LocalMux I__4694 (
            .O(N__23994),
            .I(N__23982));
    InMux I__4693 (
            .O(N__23993),
            .I(N__23979));
    CascadeMux I__4692 (
            .O(N__23992),
            .I(N__23975));
    LocalMux I__4691 (
            .O(N__23989),
            .I(N__23971));
    LocalMux I__4690 (
            .O(N__23986),
            .I(N__23968));
    InMux I__4689 (
            .O(N__23985),
            .I(N__23965));
    Span4Mux_v I__4688 (
            .O(N__23982),
            .I(N__23960));
    LocalMux I__4687 (
            .O(N__23979),
            .I(N__23960));
    InMux I__4686 (
            .O(N__23978),
            .I(N__23957));
    InMux I__4685 (
            .O(N__23975),
            .I(N__23952));
    InMux I__4684 (
            .O(N__23974),
            .I(N__23952));
    Odrv12 I__4683 (
            .O(N__23971),
            .I(cmd_16));
    Odrv4 I__4682 (
            .O(N__23968),
            .I(cmd_16));
    LocalMux I__4681 (
            .O(N__23965),
            .I(cmd_16));
    Odrv4 I__4680 (
            .O(N__23960),
            .I(cmd_16));
    LocalMux I__4679 (
            .O(N__23957),
            .I(cmd_16));
    LocalMux I__4678 (
            .O(N__23952),
            .I(cmd_16));
    CascadeMux I__4677 (
            .O(N__23939),
            .I(N__23936));
    InMux I__4676 (
            .O(N__23936),
            .I(N__23933));
    LocalMux I__4675 (
            .O(N__23933),
            .I(N__23929));
    InMux I__4674 (
            .O(N__23932),
            .I(N__23926));
    Odrv4 I__4673 (
            .O(N__23929),
            .I(configRegister_15_adj_1345));
    LocalMux I__4672 (
            .O(N__23926),
            .I(configRegister_15_adj_1345));
    CascadeMux I__4671 (
            .O(N__23921),
            .I(N__23913));
    InMux I__4670 (
            .O(N__23920),
            .I(N__23904));
    InMux I__4669 (
            .O(N__23919),
            .I(N__23904));
    InMux I__4668 (
            .O(N__23918),
            .I(N__23904));
    InMux I__4667 (
            .O(N__23917),
            .I(N__23901));
    InMux I__4666 (
            .O(N__23916),
            .I(N__23892));
    InMux I__4665 (
            .O(N__23913),
            .I(N__23892));
    InMux I__4664 (
            .O(N__23912),
            .I(N__23892));
    InMux I__4663 (
            .O(N__23911),
            .I(N__23892));
    LocalMux I__4662 (
            .O(N__23904),
            .I(N__23885));
    LocalMux I__4661 (
            .O(N__23901),
            .I(N__23885));
    LocalMux I__4660 (
            .O(N__23892),
            .I(N__23885));
    Odrv12 I__4659 (
            .O(N__23885),
            .I(wrtrigmask_3));
    InMux I__4658 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__4657 (
            .O(N__23879),
            .I(N__23875));
    InMux I__4656 (
            .O(N__23878),
            .I(N__23872));
    Odrv4 I__4655 (
            .O(N__23875),
            .I(configRegister_12_adj_1388));
    LocalMux I__4654 (
            .O(N__23872),
            .I(configRegister_12_adj_1388));
    InMux I__4653 (
            .O(N__23867),
            .I(N__23864));
    LocalMux I__4652 (
            .O(N__23864),
            .I(N__23860));
    InMux I__4651 (
            .O(N__23863),
            .I(N__23857));
    Odrv4 I__4650 (
            .O(N__23860),
            .I(configRegister_5_adj_1355));
    LocalMux I__4649 (
            .O(N__23857),
            .I(configRegister_5_adj_1355));
    InMux I__4648 (
            .O(N__23852),
            .I(N__23849));
    LocalMux I__4647 (
            .O(N__23849),
            .I(N__23845));
    InMux I__4646 (
            .O(N__23848),
            .I(N__23842));
    Odrv12 I__4645 (
            .O(N__23845),
            .I(configRegister_14_adj_1346));
    LocalMux I__4644 (
            .O(N__23842),
            .I(configRegister_14_adj_1346));
    InMux I__4643 (
            .O(N__23837),
            .I(N__23834));
    LocalMux I__4642 (
            .O(N__23834),
            .I(N__23830));
    InMux I__4641 (
            .O(N__23833),
            .I(N__23827));
    Odrv4 I__4640 (
            .O(N__23830),
            .I(configRegister_9_adj_1351));
    LocalMux I__4639 (
            .O(N__23827),
            .I(configRegister_9_adj_1351));
    InMux I__4638 (
            .O(N__23822),
            .I(N__23818));
    InMux I__4637 (
            .O(N__23821),
            .I(N__23815));
    LocalMux I__4636 (
            .O(N__23818),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12 ));
    LocalMux I__4635 (
            .O(N__23815),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12 ));
    InMux I__4634 (
            .O(N__23810),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7910 ));
    CascadeMux I__4633 (
            .O(N__23807),
            .I(N__23804));
    InMux I__4632 (
            .O(N__23804),
            .I(N__23800));
    InMux I__4631 (
            .O(N__23803),
            .I(N__23797));
    LocalMux I__4630 (
            .O(N__23800),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13 ));
    LocalMux I__4629 (
            .O(N__23797),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13 ));
    InMux I__4628 (
            .O(N__23792),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7911 ));
    InMux I__4627 (
            .O(N__23789),
            .I(N__23785));
    InMux I__4626 (
            .O(N__23788),
            .I(N__23782));
    LocalMux I__4625 (
            .O(N__23785),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14 ));
    LocalMux I__4624 (
            .O(N__23782),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14 ));
    InMux I__4623 (
            .O(N__23777),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7912 ));
    CascadeMux I__4622 (
            .O(N__23774),
            .I(N__23766));
    CascadeMux I__4621 (
            .O(N__23773),
            .I(N__23762));
    CascadeMux I__4620 (
            .O(N__23772),
            .I(N__23758));
    CascadeMux I__4619 (
            .O(N__23771),
            .I(N__23754));
    CascadeMux I__4618 (
            .O(N__23770),
            .I(N__23748));
    InMux I__4617 (
            .O(N__23769),
            .I(N__23745));
    InMux I__4616 (
            .O(N__23766),
            .I(N__23730));
    InMux I__4615 (
            .O(N__23765),
            .I(N__23730));
    InMux I__4614 (
            .O(N__23762),
            .I(N__23730));
    InMux I__4613 (
            .O(N__23761),
            .I(N__23730));
    InMux I__4612 (
            .O(N__23758),
            .I(N__23730));
    InMux I__4611 (
            .O(N__23757),
            .I(N__23730));
    InMux I__4610 (
            .O(N__23754),
            .I(N__23730));
    CascadeMux I__4609 (
            .O(N__23753),
            .I(N__23726));
    CascadeMux I__4608 (
            .O(N__23752),
            .I(N__23722));
    CascadeMux I__4607 (
            .O(N__23751),
            .I(N__23718));
    InMux I__4606 (
            .O(N__23748),
            .I(N__23715));
    LocalMux I__4605 (
            .O(N__23745),
            .I(N__23710));
    LocalMux I__4604 (
            .O(N__23730),
            .I(N__23710));
    InMux I__4603 (
            .O(N__23729),
            .I(N__23697));
    InMux I__4602 (
            .O(N__23726),
            .I(N__23697));
    InMux I__4601 (
            .O(N__23725),
            .I(N__23697));
    InMux I__4600 (
            .O(N__23722),
            .I(N__23697));
    InMux I__4599 (
            .O(N__23721),
            .I(N__23697));
    InMux I__4598 (
            .O(N__23718),
            .I(N__23697));
    LocalMux I__4597 (
            .O(N__23715),
            .I(N__23694));
    Odrv4 I__4596 (
            .O(N__23710),
            .I(\Inst_core.n1639 ));
    LocalMux I__4595 (
            .O(N__23697),
            .I(\Inst_core.n1639 ));
    Odrv4 I__4594 (
            .O(N__23694),
            .I(\Inst_core.n1639 ));
    InMux I__4593 (
            .O(N__23687),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7913 ));
    CascadeMux I__4592 (
            .O(N__23684),
            .I(N__23680));
    InMux I__4591 (
            .O(N__23683),
            .I(N__23677));
    InMux I__4590 (
            .O(N__23680),
            .I(N__23674));
    LocalMux I__4589 (
            .O(N__23677),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15 ));
    LocalMux I__4588 (
            .O(N__23674),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15 ));
    CEMux I__4587 (
            .O(N__23669),
            .I(N__23665));
    CEMux I__4586 (
            .O(N__23668),
            .I(N__23662));
    LocalMux I__4585 (
            .O(N__23665),
            .I(N__23659));
    LocalMux I__4584 (
            .O(N__23662),
            .I(N__23656));
    Span4Mux_s3_v I__4583 (
            .O(N__23659),
            .I(N__23653));
    Span4Mux_v I__4582 (
            .O(N__23656),
            .I(N__23650));
    Span4Mux_s3_h I__4581 (
            .O(N__23653),
            .I(N__23647));
    Odrv4 I__4580 (
            .O(N__23650),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4114 ));
    Odrv4 I__4579 (
            .O(N__23647),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4114 ));
    InMux I__4578 (
            .O(N__23642),
            .I(N__23637));
    InMux I__4577 (
            .O(N__23641),
            .I(N__23634));
    InMux I__4576 (
            .O(N__23640),
            .I(N__23631));
    LocalMux I__4575 (
            .O(N__23637),
            .I(N__23628));
    LocalMux I__4574 (
            .O(N__23634),
            .I(N__23625));
    LocalMux I__4573 (
            .O(N__23631),
            .I(\Inst_core.configRegister_27 ));
    Odrv4 I__4572 (
            .O(N__23628),
            .I(\Inst_core.configRegister_27 ));
    Odrv12 I__4571 (
            .O(N__23625),
            .I(\Inst_core.configRegister_27 ));
    InMux I__4570 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__4569 (
            .O(N__23615),
            .I(N__23611));
    InMux I__4568 (
            .O(N__23614),
            .I(N__23608));
    Odrv12 I__4567 (
            .O(N__23611),
            .I(configRegister_7_adj_1353));
    LocalMux I__4566 (
            .O(N__23608),
            .I(configRegister_7_adj_1353));
    InMux I__4565 (
            .O(N__23603),
            .I(N__23599));
    InMux I__4564 (
            .O(N__23602),
            .I(N__23596));
    LocalMux I__4563 (
            .O(N__23599),
            .I(configRegister_11_adj_1349));
    LocalMux I__4562 (
            .O(N__23596),
            .I(configRegister_11_adj_1349));
    CascadeMux I__4561 (
            .O(N__23591),
            .I(N__23588));
    InMux I__4560 (
            .O(N__23588),
            .I(N__23584));
    InMux I__4559 (
            .O(N__23587),
            .I(N__23581));
    LocalMux I__4558 (
            .O(N__23584),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3 ));
    LocalMux I__4557 (
            .O(N__23581),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3 ));
    InMux I__4556 (
            .O(N__23576),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7901 ));
    CascadeMux I__4555 (
            .O(N__23573),
            .I(N__23570));
    InMux I__4554 (
            .O(N__23570),
            .I(N__23566));
    InMux I__4553 (
            .O(N__23569),
            .I(N__23563));
    LocalMux I__4552 (
            .O(N__23566),
            .I(N__23560));
    LocalMux I__4551 (
            .O(N__23563),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4 ));
    Odrv4 I__4550 (
            .O(N__23560),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4 ));
    InMux I__4549 (
            .O(N__23555),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7902 ));
    CascadeMux I__4548 (
            .O(N__23552),
            .I(N__23548));
    CascadeMux I__4547 (
            .O(N__23551),
            .I(N__23545));
    InMux I__4546 (
            .O(N__23548),
            .I(N__23542));
    InMux I__4545 (
            .O(N__23545),
            .I(N__23539));
    LocalMux I__4544 (
            .O(N__23542),
            .I(N__23536));
    LocalMux I__4543 (
            .O(N__23539),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5 ));
    Odrv4 I__4542 (
            .O(N__23536),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5 ));
    InMux I__4541 (
            .O(N__23531),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7903 ));
    InMux I__4540 (
            .O(N__23528),
            .I(N__23524));
    InMux I__4539 (
            .O(N__23527),
            .I(N__23521));
    LocalMux I__4538 (
            .O(N__23524),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6 ));
    LocalMux I__4537 (
            .O(N__23521),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6 ));
    InMux I__4536 (
            .O(N__23516),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7904 ));
    CascadeMux I__4535 (
            .O(N__23513),
            .I(N__23509));
    CascadeMux I__4534 (
            .O(N__23512),
            .I(N__23506));
    InMux I__4533 (
            .O(N__23509),
            .I(N__23503));
    InMux I__4532 (
            .O(N__23506),
            .I(N__23500));
    LocalMux I__4531 (
            .O(N__23503),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7 ));
    LocalMux I__4530 (
            .O(N__23500),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7 ));
    InMux I__4529 (
            .O(N__23495),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7905 ));
    InMux I__4528 (
            .O(N__23492),
            .I(N__23488));
    InMux I__4527 (
            .O(N__23491),
            .I(N__23485));
    LocalMux I__4526 (
            .O(N__23488),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8 ));
    LocalMux I__4525 (
            .O(N__23485),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8 ));
    InMux I__4524 (
            .O(N__23480),
            .I(bfn_8_3_0_));
    CascadeMux I__4523 (
            .O(N__23477),
            .I(N__23474));
    InMux I__4522 (
            .O(N__23474),
            .I(N__23470));
    InMux I__4521 (
            .O(N__23473),
            .I(N__23467));
    LocalMux I__4520 (
            .O(N__23470),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9 ));
    LocalMux I__4519 (
            .O(N__23467),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9 ));
    InMux I__4518 (
            .O(N__23462),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7907 ));
    InMux I__4517 (
            .O(N__23459),
            .I(N__23455));
    InMux I__4516 (
            .O(N__23458),
            .I(N__23452));
    LocalMux I__4515 (
            .O(N__23455),
            .I(configRegister_10_adj_1350));
    LocalMux I__4514 (
            .O(N__23452),
            .I(configRegister_10_adj_1350));
    InMux I__4513 (
            .O(N__23447),
            .I(N__23443));
    InMux I__4512 (
            .O(N__23446),
            .I(N__23440));
    LocalMux I__4511 (
            .O(N__23443),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10 ));
    LocalMux I__4510 (
            .O(N__23440),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10 ));
    InMux I__4509 (
            .O(N__23435),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7908 ));
    CascadeMux I__4508 (
            .O(N__23432),
            .I(N__23429));
    InMux I__4507 (
            .O(N__23429),
            .I(N__23425));
    InMux I__4506 (
            .O(N__23428),
            .I(N__23422));
    LocalMux I__4505 (
            .O(N__23425),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11 ));
    LocalMux I__4504 (
            .O(N__23422),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11 ));
    InMux I__4503 (
            .O(N__23417),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7909 ));
    CascadeMux I__4502 (
            .O(N__23414),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n8808_cascade_ ));
    SRMux I__4501 (
            .O(N__23411),
            .I(N__23408));
    LocalMux I__4500 (
            .O(N__23408),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n3 ));
    CascadeMux I__4499 (
            .O(N__23405),
            .I(\Inst_core.n1639_cascade_ ));
    InMux I__4498 (
            .O(N__23402),
            .I(N__23399));
    LocalMux I__4497 (
            .O(N__23399),
            .I(\Inst_core.n9054 ));
    CascadeMux I__4496 (
            .O(N__23396),
            .I(N__23393));
    InMux I__4495 (
            .O(N__23393),
            .I(N__23389));
    InMux I__4494 (
            .O(N__23392),
            .I(N__23386));
    LocalMux I__4493 (
            .O(N__23389),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0 ));
    LocalMux I__4492 (
            .O(N__23386),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0 ));
    InMux I__4491 (
            .O(N__23381),
            .I(bfn_8_2_0_));
    InMux I__4490 (
            .O(N__23378),
            .I(N__23375));
    LocalMux I__4489 (
            .O(N__23375),
            .I(N__23371));
    InMux I__4488 (
            .O(N__23374),
            .I(N__23368));
    Odrv4 I__4487 (
            .O(N__23371),
            .I(configRegister_1_adj_1359));
    LocalMux I__4486 (
            .O(N__23368),
            .I(configRegister_1_adj_1359));
    InMux I__4485 (
            .O(N__23363),
            .I(N__23359));
    InMux I__4484 (
            .O(N__23362),
            .I(N__23356));
    LocalMux I__4483 (
            .O(N__23359),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1 ));
    LocalMux I__4482 (
            .O(N__23356),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1 ));
    InMux I__4481 (
            .O(N__23351),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7899 ));
    InMux I__4480 (
            .O(N__23348),
            .I(N__23345));
    LocalMux I__4479 (
            .O(N__23345),
            .I(N__23341));
    InMux I__4478 (
            .O(N__23344),
            .I(N__23338));
    Odrv4 I__4477 (
            .O(N__23341),
            .I(configRegister_2_adj_1358));
    LocalMux I__4476 (
            .O(N__23338),
            .I(configRegister_2_adj_1358));
    InMux I__4475 (
            .O(N__23333),
            .I(N__23329));
    InMux I__4474 (
            .O(N__23332),
            .I(N__23326));
    LocalMux I__4473 (
            .O(N__23329),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2 ));
    LocalMux I__4472 (
            .O(N__23326),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2 ));
    InMux I__4471 (
            .O(N__23321),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7900 ));
    InMux I__4470 (
            .O(N__23318),
            .I(N__23315));
    LocalMux I__4469 (
            .O(N__23315),
            .I(N__23311));
    InMux I__4468 (
            .O(N__23314),
            .I(N__23308));
    Odrv12 I__4467 (
            .O(N__23311),
            .I(configRegister_3_adj_1357));
    LocalMux I__4466 (
            .O(N__23308),
            .I(configRegister_3_adj_1357));
    InMux I__4465 (
            .O(N__23303),
            .I(N__23299));
    InMux I__4464 (
            .O(N__23302),
            .I(N__23296));
    LocalMux I__4463 (
            .O(N__23299),
            .I(N__23293));
    LocalMux I__4462 (
            .O(N__23296),
            .I(N__23290));
    Span4Mux_h I__4461 (
            .O(N__23293),
            .I(N__23287));
    Span12Mux_s11_h I__4460 (
            .O(N__23290),
            .I(N__23284));
    Span4Mux_h I__4459 (
            .O(N__23287),
            .I(N__23281));
    Odrv12 I__4458 (
            .O(N__23284),
            .I(input_c_1));
    Odrv4 I__4457 (
            .O(N__23281),
            .I(input_c_1));
    InMux I__4456 (
            .O(N__23276),
            .I(N__23272));
    InMux I__4455 (
            .O(N__23275),
            .I(N__23269));
    LocalMux I__4454 (
            .O(N__23272),
            .I(N__23266));
    LocalMux I__4453 (
            .O(N__23269),
            .I(\Inst_core.Inst_sync.synchronizedInput180_1 ));
    Odrv4 I__4452 (
            .O(N__23266),
            .I(\Inst_core.Inst_sync.synchronizedInput180_1 ));
    InMux I__4451 (
            .O(N__23261),
            .I(N__23258));
    LocalMux I__4450 (
            .O(N__23258),
            .I(N__23254));
    InMux I__4449 (
            .O(N__23257),
            .I(N__23251));
    Span4Mux_v I__4448 (
            .O(N__23254),
            .I(N__23246));
    LocalMux I__4447 (
            .O(N__23251),
            .I(N__23246));
    Span4Mux_h I__4446 (
            .O(N__23246),
            .I(N__23243));
    Odrv4 I__4445 (
            .O(N__23243),
            .I(input_c_2));
    InMux I__4444 (
            .O(N__23240),
            .I(N__23234));
    InMux I__4443 (
            .O(N__23239),
            .I(N__23234));
    LocalMux I__4442 (
            .O(N__23234),
            .I(N__23231));
    Odrv4 I__4441 (
            .O(N__23231),
            .I(\Inst_core.Inst_sync.synchronizedInput180_2 ));
    InMux I__4440 (
            .O(N__23228),
            .I(N__23224));
    InMux I__4439 (
            .O(N__23227),
            .I(N__23221));
    LocalMux I__4438 (
            .O(N__23224),
            .I(N__23218));
    LocalMux I__4437 (
            .O(N__23221),
            .I(N__23215));
    Span4Mux_h I__4436 (
            .O(N__23218),
            .I(N__23212));
    Span4Mux_h I__4435 (
            .O(N__23215),
            .I(N__23209));
    Odrv4 I__4434 (
            .O(N__23212),
            .I(input_c_3));
    Odrv4 I__4433 (
            .O(N__23209),
            .I(input_c_3));
    InMux I__4432 (
            .O(N__23204),
            .I(N__23200));
    InMux I__4431 (
            .O(N__23203),
            .I(N__23197));
    LocalMux I__4430 (
            .O(N__23200),
            .I(N__23194));
    LocalMux I__4429 (
            .O(N__23197),
            .I(\Inst_core.Inst_sync.synchronizedInput180_3 ));
    Odrv4 I__4428 (
            .O(N__23194),
            .I(\Inst_core.Inst_sync.synchronizedInput180_3 ));
    InMux I__4427 (
            .O(N__23189),
            .I(N__23185));
    InMux I__4426 (
            .O(N__23188),
            .I(N__23182));
    LocalMux I__4425 (
            .O(N__23185),
            .I(N__23179));
    LocalMux I__4424 (
            .O(N__23182),
            .I(N__23176));
    IoSpan4Mux I__4423 (
            .O(N__23179),
            .I(N__23173));
    Span4Mux_h I__4422 (
            .O(N__23176),
            .I(N__23170));
    Odrv4 I__4421 (
            .O(N__23173),
            .I(input_c_6));
    Odrv4 I__4420 (
            .O(N__23170),
            .I(input_c_6));
    InMux I__4419 (
            .O(N__23165),
            .I(N__23162));
    LocalMux I__4418 (
            .O(N__23162),
            .I(N__23158));
    InMux I__4417 (
            .O(N__23161),
            .I(N__23155));
    Odrv4 I__4416 (
            .O(N__23158),
            .I(\Inst_core.Inst_sync.synchronizedInput180_6 ));
    LocalMux I__4415 (
            .O(N__23155),
            .I(\Inst_core.Inst_sync.synchronizedInput180_6 ));
    InMux I__4414 (
            .O(N__23150),
            .I(N__23146));
    InMux I__4413 (
            .O(N__23149),
            .I(N__23143));
    LocalMux I__4412 (
            .O(N__23146),
            .I(N__23140));
    LocalMux I__4411 (
            .O(N__23143),
            .I(N__23137));
    IoSpan4Mux I__4410 (
            .O(N__23140),
            .I(N__23134));
    Span4Mux_h I__4409 (
            .O(N__23137),
            .I(N__23131));
    Odrv4 I__4408 (
            .O(N__23134),
            .I(input_c_5));
    Odrv4 I__4407 (
            .O(N__23131),
            .I(input_c_5));
    InMux I__4406 (
            .O(N__23126),
            .I(N__23123));
    LocalMux I__4405 (
            .O(N__23123),
            .I(N__23119));
    InMux I__4404 (
            .O(N__23122),
            .I(N__23116));
    Odrv4 I__4403 (
            .O(N__23119),
            .I(\Inst_core.Inst_sync.synchronizedInput180_5 ));
    LocalMux I__4402 (
            .O(N__23116),
            .I(\Inst_core.Inst_sync.synchronizedInput180_5 ));
    InMux I__4401 (
            .O(N__23111),
            .I(N__23107));
    InMux I__4400 (
            .O(N__23110),
            .I(N__23104));
    LocalMux I__4399 (
            .O(N__23107),
            .I(\Inst_core.Inst_sync.synchronizedInput180_7 ));
    LocalMux I__4398 (
            .O(N__23104),
            .I(\Inst_core.Inst_sync.synchronizedInput180_7 ));
    CascadeMux I__4397 (
            .O(N__23099),
            .I(\Inst_core.n8518_cascade_ ));
    InMux I__4396 (
            .O(N__23096),
            .I(N__23093));
    LocalMux I__4395 (
            .O(N__23093),
            .I(N__23090));
    Span12Mux_s10_v I__4394 (
            .O(N__23090),
            .I(N__23086));
    InMux I__4393 (
            .O(N__23089),
            .I(N__23083));
    Odrv12 I__4392 (
            .O(N__23086),
            .I(valueRegister_7_adj_1289));
    LocalMux I__4391 (
            .O(N__23083),
            .I(valueRegister_7_adj_1289));
    CascadeMux I__4390 (
            .O(N__23078),
            .I(N__23075));
    InMux I__4389 (
            .O(N__23075),
            .I(N__23072));
    LocalMux I__4388 (
            .O(N__23072),
            .I(N__23069));
    Span4Mux_s2_v I__4387 (
            .O(N__23069),
            .I(N__23066));
    Span4Mux_h I__4386 (
            .O(N__23066),
            .I(N__23063));
    Span4Mux_v I__4385 (
            .O(N__23063),
            .I(N__23060));
    Span4Mux_v I__4384 (
            .O(N__23060),
            .I(N__23057));
    Odrv4 I__4383 (
            .O(N__23057),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_7 ));
    InMux I__4382 (
            .O(N__23054),
            .I(N__23050));
    InMux I__4381 (
            .O(N__23053),
            .I(N__23047));
    LocalMux I__4380 (
            .O(N__23050),
            .I(N__23043));
    LocalMux I__4379 (
            .O(N__23047),
            .I(N__23040));
    InMux I__4378 (
            .O(N__23046),
            .I(N__23033));
    Span4Mux_h I__4377 (
            .O(N__23043),
            .I(N__23030));
    Span4Mux_h I__4376 (
            .O(N__23040),
            .I(N__23027));
    InMux I__4375 (
            .O(N__23039),
            .I(N__23022));
    InMux I__4374 (
            .O(N__23038),
            .I(N__23019));
    InMux I__4373 (
            .O(N__23037),
            .I(N__23015));
    InMux I__4372 (
            .O(N__23036),
            .I(N__23012));
    LocalMux I__4371 (
            .O(N__23033),
            .I(N__23009));
    Span4Mux_v I__4370 (
            .O(N__23030),
            .I(N__23006));
    Sp12to4 I__4369 (
            .O(N__23027),
            .I(N__23003));
    InMux I__4368 (
            .O(N__23026),
            .I(N__23000));
    InMux I__4367 (
            .O(N__23025),
            .I(N__22997));
    LocalMux I__4366 (
            .O(N__23022),
            .I(N__22994));
    LocalMux I__4365 (
            .O(N__23019),
            .I(N__22991));
    InMux I__4364 (
            .O(N__23018),
            .I(N__22988));
    LocalMux I__4363 (
            .O(N__23015),
            .I(N__22983));
    LocalMux I__4362 (
            .O(N__23012),
            .I(N__22983));
    Span4Mux_v I__4361 (
            .O(N__23009),
            .I(N__22980));
    Span4Mux_v I__4360 (
            .O(N__23006),
            .I(N__22977));
    Span12Mux_s5_v I__4359 (
            .O(N__23003),
            .I(N__22970));
    LocalMux I__4358 (
            .O(N__23000),
            .I(N__22970));
    LocalMux I__4357 (
            .O(N__22997),
            .I(N__22970));
    Span4Mux_v I__4356 (
            .O(N__22994),
            .I(N__22965));
    Span4Mux_h I__4355 (
            .O(N__22991),
            .I(N__22965));
    LocalMux I__4354 (
            .O(N__22988),
            .I(memoryOut_7));
    Odrv12 I__4353 (
            .O(N__22983),
            .I(memoryOut_7));
    Odrv4 I__4352 (
            .O(N__22980),
            .I(memoryOut_7));
    Odrv4 I__4351 (
            .O(N__22977),
            .I(memoryOut_7));
    Odrv12 I__4350 (
            .O(N__22970),
            .I(memoryOut_7));
    Odrv4 I__4349 (
            .O(N__22965),
            .I(memoryOut_7));
    InMux I__4348 (
            .O(N__22952),
            .I(N__22948));
    InMux I__4347 (
            .O(N__22951),
            .I(N__22945));
    LocalMux I__4346 (
            .O(N__22948),
            .I(N__22942));
    LocalMux I__4345 (
            .O(N__22945),
            .I(N__22939));
    Span4Mux_v I__4344 (
            .O(N__22942),
            .I(N__22936));
    Odrv12 I__4343 (
            .O(N__22939),
            .I(\Inst_core.Inst_sync.demuxedInput_7 ));
    Odrv4 I__4342 (
            .O(N__22936),
            .I(\Inst_core.Inst_sync.demuxedInput_7 ));
    InMux I__4341 (
            .O(N__22931),
            .I(N__22927));
    InMux I__4340 (
            .O(N__22930),
            .I(N__22924));
    LocalMux I__4339 (
            .O(N__22927),
            .I(N__22921));
    LocalMux I__4338 (
            .O(N__22924),
            .I(N__22917));
    Span4Mux_v I__4337 (
            .O(N__22921),
            .I(N__22914));
    InMux I__4336 (
            .O(N__22920),
            .I(N__22911));
    Span4Mux_h I__4335 (
            .O(N__22917),
            .I(N__22908));
    Span4Mux_h I__4334 (
            .O(N__22914),
            .I(N__22905));
    LocalMux I__4333 (
            .O(N__22911),
            .I(N__22902));
    Odrv4 I__4332 (
            .O(N__22908),
            .I(\Inst_core.Inst_sync.demuxedInput_2 ));
    Odrv4 I__4331 (
            .O(N__22905),
            .I(\Inst_core.Inst_sync.demuxedInput_2 ));
    Odrv4 I__4330 (
            .O(N__22902),
            .I(\Inst_core.Inst_sync.demuxedInput_2 ));
    InMux I__4329 (
            .O(N__22895),
            .I(N__22891));
    InMux I__4328 (
            .O(N__22894),
            .I(N__22888));
    LocalMux I__4327 (
            .O(N__22891),
            .I(N__22885));
    LocalMux I__4326 (
            .O(N__22888),
            .I(N__22882));
    Span4Mux_h I__4325 (
            .O(N__22885),
            .I(N__22879));
    Odrv4 I__4324 (
            .O(N__22882),
            .I(\Inst_core.Inst_sync.demuxedInput_5 ));
    Odrv4 I__4323 (
            .O(N__22879),
            .I(\Inst_core.Inst_sync.demuxedInput_5 ));
    InMux I__4322 (
            .O(N__22874),
            .I(N__22871));
    LocalMux I__4321 (
            .O(N__22871),
            .I(N__22868));
    Odrv4 I__4320 (
            .O(N__22868),
            .I(\Inst_core.Inst_sync.n9117 ));
    InMux I__4319 (
            .O(N__22865),
            .I(N__22861));
    InMux I__4318 (
            .O(N__22864),
            .I(N__22858));
    LocalMux I__4317 (
            .O(N__22861),
            .I(N__22855));
    LocalMux I__4316 (
            .O(N__22858),
            .I(N__22850));
    Span4Mux_h I__4315 (
            .O(N__22855),
            .I(N__22850));
    Span4Mux_v I__4314 (
            .O(N__22850),
            .I(N__22846));
    InMux I__4313 (
            .O(N__22849),
            .I(N__22843));
    Span4Mux_v I__4312 (
            .O(N__22846),
            .I(N__22840));
    LocalMux I__4311 (
            .O(N__22843),
            .I(N__22837));
    Odrv4 I__4310 (
            .O(N__22840),
            .I(\Inst_core.Inst_sync.demuxedInput_3 ));
    Odrv4 I__4309 (
            .O(N__22837),
            .I(\Inst_core.Inst_sync.demuxedInput_3 ));
    CascadeMux I__4308 (
            .O(N__22832),
            .I(N__22829));
    InMux I__4307 (
            .O(N__22829),
            .I(N__22824));
    InMux I__4306 (
            .O(N__22828),
            .I(N__22821));
    InMux I__4305 (
            .O(N__22827),
            .I(N__22818));
    LocalMux I__4304 (
            .O(N__22824),
            .I(N__22815));
    LocalMux I__4303 (
            .O(N__22821),
            .I(\Inst_core.Inst_sync.synchronizedInput_5 ));
    LocalMux I__4302 (
            .O(N__22818),
            .I(\Inst_core.Inst_sync.synchronizedInput_5 ));
    Odrv4 I__4301 (
            .O(N__22815),
            .I(\Inst_core.Inst_sync.synchronizedInput_5 ));
    InMux I__4300 (
            .O(N__22808),
            .I(N__22796));
    InMux I__4299 (
            .O(N__22807),
            .I(N__22796));
    InMux I__4298 (
            .O(N__22806),
            .I(N__22791));
    InMux I__4297 (
            .O(N__22805),
            .I(N__22791));
    InMux I__4296 (
            .O(N__22804),
            .I(N__22788));
    InMux I__4295 (
            .O(N__22803),
            .I(N__22785));
    InMux I__4294 (
            .O(N__22802),
            .I(N__22780));
    InMux I__4293 (
            .O(N__22801),
            .I(N__22780));
    LocalMux I__4292 (
            .O(N__22796),
            .I(N__22775));
    LocalMux I__4291 (
            .O(N__22791),
            .I(N__22775));
    LocalMux I__4290 (
            .O(N__22788),
            .I(\Inst_core.Inst_sync.n2566 ));
    LocalMux I__4289 (
            .O(N__22785),
            .I(\Inst_core.Inst_sync.n2566 ));
    LocalMux I__4288 (
            .O(N__22780),
            .I(\Inst_core.Inst_sync.n2566 ));
    Odrv4 I__4287 (
            .O(N__22775),
            .I(\Inst_core.Inst_sync.n2566 ));
    InMux I__4286 (
            .O(N__22766),
            .I(N__22754));
    InMux I__4285 (
            .O(N__22765),
            .I(N__22754));
    InMux I__4284 (
            .O(N__22764),
            .I(N__22754));
    InMux I__4283 (
            .O(N__22763),
            .I(N__22754));
    LocalMux I__4282 (
            .O(N__22754),
            .I(N__22747));
    InMux I__4281 (
            .O(N__22753),
            .I(N__22742));
    InMux I__4280 (
            .O(N__22752),
            .I(N__22742));
    InMux I__4279 (
            .O(N__22751),
            .I(N__22739));
    InMux I__4278 (
            .O(N__22750),
            .I(N__22736));
    Span4Mux_h I__4277 (
            .O(N__22747),
            .I(N__22733));
    LocalMux I__4276 (
            .O(N__22742),
            .I(N__22730));
    LocalMux I__4275 (
            .O(N__22739),
            .I(\Inst_core.Inst_sync.n2564 ));
    LocalMux I__4274 (
            .O(N__22736),
            .I(\Inst_core.Inst_sync.n2564 ));
    Odrv4 I__4273 (
            .O(N__22733),
            .I(\Inst_core.Inst_sync.n2564 ));
    Odrv4 I__4272 (
            .O(N__22730),
            .I(\Inst_core.Inst_sync.n2564 ));
    InMux I__4271 (
            .O(N__22721),
            .I(N__22718));
    LocalMux I__4270 (
            .O(N__22718),
            .I(N__22715));
    Odrv4 I__4269 (
            .O(N__22715),
            .I(\Inst_core.Inst_sync.n9129 ));
    InMux I__4268 (
            .O(N__22712),
            .I(N__22708));
    InMux I__4267 (
            .O(N__22711),
            .I(N__22704));
    LocalMux I__4266 (
            .O(N__22708),
            .I(N__22701));
    CascadeMux I__4265 (
            .O(N__22707),
            .I(N__22698));
    LocalMux I__4264 (
            .O(N__22704),
            .I(N__22693));
    Span4Mux_h I__4263 (
            .O(N__22701),
            .I(N__22693));
    InMux I__4262 (
            .O(N__22698),
            .I(N__22690));
    Odrv4 I__4261 (
            .O(N__22693),
            .I(\Inst_core.Inst_sync.synchronizedInput_6 ));
    LocalMux I__4260 (
            .O(N__22690),
            .I(\Inst_core.Inst_sync.synchronizedInput_6 ));
    InMux I__4259 (
            .O(N__22685),
            .I(N__22682));
    LocalMux I__4258 (
            .O(N__22682),
            .I(N__22678));
    InMux I__4257 (
            .O(N__22681),
            .I(N__22675));
    Span4Mux_h I__4256 (
            .O(N__22678),
            .I(N__22670));
    LocalMux I__4255 (
            .O(N__22675),
            .I(N__22670));
    Span4Mux_h I__4254 (
            .O(N__22670),
            .I(N__22667));
    IoSpan4Mux I__4253 (
            .O(N__22667),
            .I(N__22664));
    Odrv4 I__4252 (
            .O(N__22664),
            .I(input_c_0));
    InMux I__4251 (
            .O(N__22661),
            .I(N__22657));
    InMux I__4250 (
            .O(N__22660),
            .I(N__22654));
    LocalMux I__4249 (
            .O(N__22657),
            .I(N__22651));
    LocalMux I__4248 (
            .O(N__22654),
            .I(\Inst_core.Inst_sync.synchronizedInput180_0 ));
    Odrv4 I__4247 (
            .O(N__22651),
            .I(\Inst_core.Inst_sync.synchronizedInput180_0 ));
    CascadeMux I__4246 (
            .O(N__22646),
            .I(N__22643));
    InMux I__4245 (
            .O(N__22643),
            .I(N__22640));
    LocalMux I__4244 (
            .O(N__22640),
            .I(N__22637));
    Span4Mux_h I__4243 (
            .O(N__22637),
            .I(N__22633));
    InMux I__4242 (
            .O(N__22636),
            .I(N__22630));
    Span4Mux_h I__4241 (
            .O(N__22633),
            .I(N__22627));
    LocalMux I__4240 (
            .O(N__22630),
            .I(\Inst_core.Inst_sync.filteredInput_0 ));
    Odrv4 I__4239 (
            .O(N__22627),
            .I(\Inst_core.Inst_sync.filteredInput_0 ));
    InMux I__4238 (
            .O(N__22622),
            .I(N__22619));
    LocalMux I__4237 (
            .O(N__22619),
            .I(\Inst_core.Inst_sync.n2793 ));
    InMux I__4236 (
            .O(N__22616),
            .I(N__22612));
    InMux I__4235 (
            .O(N__22615),
            .I(N__22609));
    LocalMux I__4234 (
            .O(N__22612),
            .I(N__22606));
    LocalMux I__4233 (
            .O(N__22609),
            .I(flagInverted));
    Odrv12 I__4232 (
            .O(N__22606),
            .I(flagInverted));
    InMux I__4231 (
            .O(N__22601),
            .I(N__22589));
    InMux I__4230 (
            .O(N__22600),
            .I(N__22589));
    InMux I__4229 (
            .O(N__22599),
            .I(N__22589));
    InMux I__4228 (
            .O(N__22598),
            .I(N__22584));
    InMux I__4227 (
            .O(N__22597),
            .I(N__22584));
    InMux I__4226 (
            .O(N__22596),
            .I(N__22580));
    LocalMux I__4225 (
            .O(N__22589),
            .I(N__22575));
    LocalMux I__4224 (
            .O(N__22584),
            .I(N__22575));
    InMux I__4223 (
            .O(N__22583),
            .I(N__22572));
    LocalMux I__4222 (
            .O(N__22580),
            .I(N__22569));
    Span4Mux_v I__4221 (
            .O(N__22575),
            .I(N__22566));
    LocalMux I__4220 (
            .O(N__22572),
            .I(flagFilter));
    Odrv12 I__4219 (
            .O(N__22569),
            .I(flagFilter));
    Odrv4 I__4218 (
            .O(N__22566),
            .I(flagFilter));
    InMux I__4217 (
            .O(N__22559),
            .I(N__22555));
    InMux I__4216 (
            .O(N__22558),
            .I(N__22552));
    LocalMux I__4215 (
            .O(N__22555),
            .I(N__22549));
    LocalMux I__4214 (
            .O(N__22552),
            .I(N__22543));
    Span4Mux_h I__4213 (
            .O(N__22549),
            .I(N__22543));
    InMux I__4212 (
            .O(N__22548),
            .I(N__22540));
    Odrv4 I__4211 (
            .O(N__22543),
            .I(\Inst_core.Inst_sync.demuxedInput_1 ));
    LocalMux I__4210 (
            .O(N__22540),
            .I(\Inst_core.Inst_sync.demuxedInput_1 ));
    InMux I__4209 (
            .O(N__22535),
            .I(N__22532));
    LocalMux I__4208 (
            .O(N__22532),
            .I(\Inst_core.Inst_sync.n2787 ));
    InMux I__4207 (
            .O(N__22529),
            .I(N__22526));
    LocalMux I__4206 (
            .O(N__22526),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_5 ));
    CascadeMux I__4205 (
            .O(N__22523),
            .I(N__22520));
    InMux I__4204 (
            .O(N__22520),
            .I(N__22517));
    LocalMux I__4203 (
            .O(N__22517),
            .I(syncedInput_6));
    InMux I__4202 (
            .O(N__22514),
            .I(N__22511));
    LocalMux I__4201 (
            .O(N__22511),
            .I(N__22508));
    Span4Mux_v I__4200 (
            .O(N__22508),
            .I(N__22505));
    Odrv4 I__4199 (
            .O(N__22505),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_6 ));
    CascadeMux I__4198 (
            .O(N__22502),
            .I(N__22499));
    InMux I__4197 (
            .O(N__22499),
            .I(N__22496));
    LocalMux I__4196 (
            .O(N__22496),
            .I(syncedInput_3));
    CascadeMux I__4195 (
            .O(N__22493),
            .I(N__22490));
    InMux I__4194 (
            .O(N__22490),
            .I(N__22487));
    LocalMux I__4193 (
            .O(N__22487),
            .I(N__22484));
    Span4Mux_h I__4192 (
            .O(N__22484),
            .I(N__22481));
    Odrv4 I__4191 (
            .O(N__22481),
            .I(syncedInput_7));
    InMux I__4190 (
            .O(N__22478),
            .I(N__22474));
    InMux I__4189 (
            .O(N__22477),
            .I(N__22471));
    LocalMux I__4188 (
            .O(N__22474),
            .I(valueRegister_7_adj_1329));
    LocalMux I__4187 (
            .O(N__22471),
            .I(valueRegister_7_adj_1329));
    CascadeMux I__4186 (
            .O(N__22466),
            .I(N__22463));
    InMux I__4185 (
            .O(N__22463),
            .I(N__22460));
    LocalMux I__4184 (
            .O(N__22460),
            .I(N__22457));
    Span4Mux_v I__4183 (
            .O(N__22457),
            .I(N__22453));
    InMux I__4182 (
            .O(N__22456),
            .I(N__22450));
    Span4Mux_h I__4181 (
            .O(N__22453),
            .I(N__22447));
    LocalMux I__4180 (
            .O(N__22450),
            .I(\Inst_core.Inst_sync.filteredInput_1 ));
    Odrv4 I__4179 (
            .O(N__22447),
            .I(\Inst_core.Inst_sync.filteredInput_1 ));
    CascadeMux I__4178 (
            .O(N__22442),
            .I(N__22439));
    InMux I__4177 (
            .O(N__22439),
            .I(N__22436));
    LocalMux I__4176 (
            .O(N__22436),
            .I(N__22432));
    InMux I__4175 (
            .O(N__22435),
            .I(N__22429));
    Span12Mux_s7_h I__4174 (
            .O(N__22432),
            .I(N__22426));
    LocalMux I__4173 (
            .O(N__22429),
            .I(\Inst_core.Inst_sync.filteredInput_3 ));
    Odrv12 I__4172 (
            .O(N__22426),
            .I(\Inst_core.Inst_sync.filteredInput_3 ));
    InMux I__4171 (
            .O(N__22421),
            .I(N__22418));
    LocalMux I__4170 (
            .O(N__22418),
            .I(\Inst_core.Inst_sync.n2791 ));
    InMux I__4169 (
            .O(N__22415),
            .I(N__22412));
    LocalMux I__4168 (
            .O(N__22412),
            .I(N__22409));
    Span4Mux_s2_h I__4167 (
            .O(N__22409),
            .I(N__22406));
    Span4Mux_h I__4166 (
            .O(N__22406),
            .I(N__22403));
    Odrv4 I__4165 (
            .O(N__22403),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_1 ));
    SRMux I__4164 (
            .O(N__22400),
            .I(N__22397));
    LocalMux I__4163 (
            .O(N__22397),
            .I(N__22394));
    Span4Mux_v I__4162 (
            .O(N__22394),
            .I(N__22391));
    Span4Mux_h I__4161 (
            .O(N__22391),
            .I(N__22388));
    Span4Mux_h I__4160 (
            .O(N__22388),
            .I(N__22385));
    Odrv4 I__4159 (
            .O(N__22385),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4746 ));
    InMux I__4158 (
            .O(N__22382),
            .I(N__22379));
    LocalMux I__4157 (
            .O(N__22379),
            .I(N__22375));
    InMux I__4156 (
            .O(N__22378),
            .I(N__22372));
    Span4Mux_v I__4155 (
            .O(N__22375),
            .I(N__22369));
    LocalMux I__4154 (
            .O(N__22372),
            .I(fwd_15));
    Odrv4 I__4153 (
            .O(N__22369),
            .I(fwd_15));
    CascadeMux I__4152 (
            .O(N__22364),
            .I(\Inst_core.Inst_controller.n22_cascade_ ));
    InMux I__4151 (
            .O(N__22361),
            .I(N__22357));
    InMux I__4150 (
            .O(N__22360),
            .I(N__22354));
    LocalMux I__4149 (
            .O(N__22357),
            .I(fwd_6));
    LocalMux I__4148 (
            .O(N__22354),
            .I(fwd_6));
    CascadeMux I__4147 (
            .O(N__22349),
            .I(\Inst_core.Inst_controller.n4_adj_986_cascade_ ));
    InMux I__4146 (
            .O(N__22346),
            .I(N__22342));
    InMux I__4145 (
            .O(N__22345),
            .I(N__22339));
    LocalMux I__4144 (
            .O(N__22342),
            .I(fwd_5));
    LocalMux I__4143 (
            .O(N__22339),
            .I(fwd_5));
    CascadeMux I__4142 (
            .O(N__22334),
            .I(\Inst_core.Inst_controller.n4_adj_987_cascade_ ));
    InMux I__4141 (
            .O(N__22331),
            .I(N__22328));
    LocalMux I__4140 (
            .O(N__22328),
            .I(\Inst_core.Inst_controller.n8486 ));
    InMux I__4139 (
            .O(N__22325),
            .I(N__22322));
    LocalMux I__4138 (
            .O(N__22322),
            .I(N__22319));
    Span4Mux_h I__4137 (
            .O(N__22319),
            .I(N__22314));
    InMux I__4136 (
            .O(N__22318),
            .I(N__22311));
    InMux I__4135 (
            .O(N__22317),
            .I(N__22308));
    Span4Mux_v I__4134 (
            .O(N__22314),
            .I(N__22305));
    LocalMux I__4133 (
            .O(N__22311),
            .I(N__22302));
    LocalMux I__4132 (
            .O(N__22308),
            .I(\Inst_core.Inst_sync.demuxedInput_0 ));
    Odrv4 I__4131 (
            .O(N__22305),
            .I(\Inst_core.Inst_sync.demuxedInput_0 ));
    Odrv12 I__4130 (
            .O(N__22302),
            .I(\Inst_core.Inst_sync.demuxedInput_0 ));
    CascadeMux I__4129 (
            .O(N__22295),
            .I(N__22292));
    InMux I__4128 (
            .O(N__22292),
            .I(N__22286));
    InMux I__4127 (
            .O(N__22291),
            .I(N__22286));
    LocalMux I__4126 (
            .O(N__22286),
            .I(N__22282));
    InMux I__4125 (
            .O(N__22285),
            .I(N__22279));
    Span4Mux_s3_h I__4124 (
            .O(N__22282),
            .I(N__22272));
    LocalMux I__4123 (
            .O(N__22279),
            .I(N__22272));
    InMux I__4122 (
            .O(N__22278),
            .I(N__22269));
    InMux I__4121 (
            .O(N__22277),
            .I(N__22266));
    Span4Mux_h I__4120 (
            .O(N__22272),
            .I(N__22261));
    LocalMux I__4119 (
            .O(N__22269),
            .I(N__22261));
    LocalMux I__4118 (
            .O(N__22266),
            .I(N__22257));
    Span4Mux_v I__4117 (
            .O(N__22261),
            .I(N__22253));
    InMux I__4116 (
            .O(N__22260),
            .I(N__22250));
    Sp12to4 I__4115 (
            .O(N__22257),
            .I(N__22247));
    InMux I__4114 (
            .O(N__22256),
            .I(N__22244));
    Sp12to4 I__4113 (
            .O(N__22253),
            .I(N__22239));
    LocalMux I__4112 (
            .O(N__22250),
            .I(N__22239));
    Span12Mux_s11_v I__4111 (
            .O(N__22247),
            .I(N__22236));
    LocalMux I__4110 (
            .O(N__22244),
            .I(N__22231));
    Span12Mux_s8_h I__4109 (
            .O(N__22239),
            .I(N__22231));
    Odrv12 I__4108 (
            .O(N__22236),
            .I(wrFlags));
    Odrv12 I__4107 (
            .O(N__22231),
            .I(wrFlags));
    InMux I__4106 (
            .O(N__22226),
            .I(N__22220));
    InMux I__4105 (
            .O(N__22225),
            .I(N__22220));
    LocalMux I__4104 (
            .O(N__22220),
            .I(N__22213));
    InMux I__4103 (
            .O(N__22219),
            .I(N__22210));
    InMux I__4102 (
            .O(N__22218),
            .I(N__22207));
    InMux I__4101 (
            .O(N__22217),
            .I(N__22204));
    CascadeMux I__4100 (
            .O(N__22216),
            .I(N__22200));
    Span4Mux_h I__4099 (
            .O(N__22213),
            .I(N__22197));
    LocalMux I__4098 (
            .O(N__22210),
            .I(N__22194));
    LocalMux I__4097 (
            .O(N__22207),
            .I(N__22189));
    LocalMux I__4096 (
            .O(N__22204),
            .I(N__22189));
    InMux I__4095 (
            .O(N__22203),
            .I(N__22186));
    InMux I__4094 (
            .O(N__22200),
            .I(N__22183));
    Odrv4 I__4093 (
            .O(N__22197),
            .I(cmd_32));
    Odrv4 I__4092 (
            .O(N__22194),
            .I(cmd_32));
    Odrv4 I__4091 (
            .O(N__22189),
            .I(cmd_32));
    LocalMux I__4090 (
            .O(N__22186),
            .I(cmd_32));
    LocalMux I__4089 (
            .O(N__22183),
            .I(cmd_32));
    InMux I__4088 (
            .O(N__22172),
            .I(N__22168));
    InMux I__4087 (
            .O(N__22171),
            .I(N__22165));
    LocalMux I__4086 (
            .O(N__22168),
            .I(N__22162));
    LocalMux I__4085 (
            .O(N__22165),
            .I(N__22158));
    Span4Mux_s2_h I__4084 (
            .O(N__22162),
            .I(N__22155));
    InMux I__4083 (
            .O(N__22161),
            .I(N__22152));
    Span4Mux_h I__4082 (
            .O(N__22158),
            .I(N__22147));
    Span4Mux_h I__4081 (
            .O(N__22155),
            .I(N__22147));
    LocalMux I__4080 (
            .O(N__22152),
            .I(configRegister_20));
    Odrv4 I__4079 (
            .O(N__22147),
            .I(configRegister_20));
    InMux I__4078 (
            .O(N__22142),
            .I(N__22139));
    LocalMux I__4077 (
            .O(N__22139),
            .I(N__22136));
    Span4Mux_v I__4076 (
            .O(N__22136),
            .I(N__22132));
    InMux I__4075 (
            .O(N__22135),
            .I(N__22129));
    Odrv4 I__4074 (
            .O(N__22132),
            .I(valueRegister_1_adj_1295));
    LocalMux I__4073 (
            .O(N__22129),
            .I(valueRegister_1_adj_1295));
    InMux I__4072 (
            .O(N__22124),
            .I(N__22119));
    InMux I__4071 (
            .O(N__22123),
            .I(N__22114));
    InMux I__4070 (
            .O(N__22122),
            .I(N__22114));
    LocalMux I__4069 (
            .O(N__22119),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1 ));
    LocalMux I__4068 (
            .O(N__22114),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1 ));
    InMux I__4067 (
            .O(N__22109),
            .I(N__22103));
    InMux I__4066 (
            .O(N__22108),
            .I(N__22103));
    LocalMux I__4065 (
            .O(N__22103),
            .I(N__22099));
    InMux I__4064 (
            .O(N__22102),
            .I(N__22096));
    Span4Mux_h I__4063 (
            .O(N__22099),
            .I(N__22093));
    LocalMux I__4062 (
            .O(N__22096),
            .I(configRegister_22_adj_1340));
    Odrv4 I__4061 (
            .O(N__22093),
            .I(configRegister_22_adj_1340));
    CascadeMux I__4060 (
            .O(N__22088),
            .I(N__22083));
    CascadeMux I__4059 (
            .O(N__22087),
            .I(N__22080));
    InMux I__4058 (
            .O(N__22086),
            .I(N__22075));
    InMux I__4057 (
            .O(N__22083),
            .I(N__22075));
    InMux I__4056 (
            .O(N__22080),
            .I(N__22071));
    LocalMux I__4055 (
            .O(N__22075),
            .I(N__22068));
    InMux I__4054 (
            .O(N__22074),
            .I(N__22065));
    LocalMux I__4053 (
            .O(N__22071),
            .I(N__22062));
    Span4Mux_v I__4052 (
            .O(N__22068),
            .I(N__22058));
    LocalMux I__4051 (
            .O(N__22065),
            .I(N__22053));
    Span4Mux_v I__4050 (
            .O(N__22062),
            .I(N__22053));
    InMux I__4049 (
            .O(N__22061),
            .I(N__22050));
    Span4Mux_h I__4048 (
            .O(N__22058),
            .I(N__22047));
    Span4Mux_h I__4047 (
            .O(N__22053),
            .I(N__22044));
    LocalMux I__4046 (
            .O(N__22050),
            .I(configRegister_21));
    Odrv4 I__4045 (
            .O(N__22047),
            .I(configRegister_21));
    Odrv4 I__4044 (
            .O(N__22044),
            .I(configRegister_21));
    InMux I__4043 (
            .O(N__22037),
            .I(N__22031));
    InMux I__4042 (
            .O(N__22036),
            .I(N__22028));
    InMux I__4041 (
            .O(N__22035),
            .I(N__22019));
    InMux I__4040 (
            .O(N__22034),
            .I(N__22019));
    LocalMux I__4039 (
            .O(N__22031),
            .I(N__22016));
    LocalMux I__4038 (
            .O(N__22028),
            .I(N__22013));
    InMux I__4037 (
            .O(N__22027),
            .I(N__22010));
    InMux I__4036 (
            .O(N__22026),
            .I(N__22007));
    InMux I__4035 (
            .O(N__22025),
            .I(N__22004));
    InMux I__4034 (
            .O(N__22024),
            .I(N__22001));
    LocalMux I__4033 (
            .O(N__22019),
            .I(N__21998));
    Span4Mux_h I__4032 (
            .O(N__22016),
            .I(N__21995));
    Span4Mux_h I__4031 (
            .O(N__22013),
            .I(N__21992));
    LocalMux I__4030 (
            .O(N__22010),
            .I(N__21985));
    LocalMux I__4029 (
            .O(N__22007),
            .I(N__21985));
    LocalMux I__4028 (
            .O(N__22004),
            .I(N__21985));
    LocalMux I__4027 (
            .O(N__22001),
            .I(N__21982));
    Span4Mux_h I__4026 (
            .O(N__21998),
            .I(N__21979));
    Span4Mux_s3_h I__4025 (
            .O(N__21995),
            .I(N__21976));
    Span4Mux_v I__4024 (
            .O(N__21992),
            .I(N__21971));
    Span4Mux_v I__4023 (
            .O(N__21985),
            .I(N__21971));
    Span12Mux_s8_h I__4022 (
            .O(N__21982),
            .I(N__21964));
    Sp12to4 I__4021 (
            .O(N__21979),
            .I(N__21964));
    Sp12to4 I__4020 (
            .O(N__21976),
            .I(N__21964));
    Odrv4 I__4019 (
            .O(N__21971),
            .I(wrtrigmask_1));
    Odrv12 I__4018 (
            .O(N__21964),
            .I(wrtrigmask_1));
    CascadeMux I__4017 (
            .O(N__21959),
            .I(N__21953));
    InMux I__4016 (
            .O(N__21958),
            .I(N__21943));
    InMux I__4015 (
            .O(N__21957),
            .I(N__21943));
    InMux I__4014 (
            .O(N__21956),
            .I(N__21943));
    InMux I__4013 (
            .O(N__21953),
            .I(N__21943));
    InMux I__4012 (
            .O(N__21952),
            .I(N__21940));
    LocalMux I__4011 (
            .O(N__21943),
            .I(N__21937));
    LocalMux I__4010 (
            .O(N__21940),
            .I(configRegister_21_adj_1341));
    Odrv4 I__4009 (
            .O(N__21937),
            .I(configRegister_21_adj_1341));
    InMux I__4008 (
            .O(N__21932),
            .I(N__21926));
    InMux I__4007 (
            .O(N__21931),
            .I(N__21926));
    LocalMux I__4006 (
            .O(N__21926),
            .I(N__21922));
    InMux I__4005 (
            .O(N__21925),
            .I(N__21919));
    Span4Mux_v I__4004 (
            .O(N__21922),
            .I(N__21916));
    LocalMux I__4003 (
            .O(N__21919),
            .I(configRegister_22_adj_1380));
    Odrv4 I__4002 (
            .O(N__21916),
            .I(configRegister_22_adj_1380));
    InMux I__4001 (
            .O(N__21911),
            .I(N__21905));
    InMux I__4000 (
            .O(N__21910),
            .I(N__21905));
    LocalMux I__3999 (
            .O(N__21905),
            .I(N__21901));
    InMux I__3998 (
            .O(N__21904),
            .I(N__21898));
    Span4Mux_h I__3997 (
            .O(N__21901),
            .I(N__21895));
    LocalMux I__3996 (
            .O(N__21898),
            .I(configRegister_23));
    Odrv4 I__3995 (
            .O(N__21895),
            .I(configRegister_23));
    InMux I__3994 (
            .O(N__21890),
            .I(N__21881));
    InMux I__3993 (
            .O(N__21889),
            .I(N__21878));
    InMux I__3992 (
            .O(N__21888),
            .I(N__21875));
    InMux I__3991 (
            .O(N__21887),
            .I(N__21866));
    InMux I__3990 (
            .O(N__21886),
            .I(N__21866));
    InMux I__3989 (
            .O(N__21885),
            .I(N__21866));
    InMux I__3988 (
            .O(N__21884),
            .I(N__21866));
    LocalMux I__3987 (
            .O(N__21881),
            .I(N__21862));
    LocalMux I__3986 (
            .O(N__21878),
            .I(N__21859));
    LocalMux I__3985 (
            .O(N__21875),
            .I(N__21856));
    LocalMux I__3984 (
            .O(N__21866),
            .I(N__21853));
    InMux I__3983 (
            .O(N__21865),
            .I(N__21850));
    Span4Mux_h I__3982 (
            .O(N__21862),
            .I(N__21847));
    Span4Mux_s3_h I__3981 (
            .O(N__21859),
            .I(N__21842));
    Span4Mux_h I__3980 (
            .O(N__21856),
            .I(N__21842));
    Span4Mux_v I__3979 (
            .O(N__21853),
            .I(N__21837));
    LocalMux I__3978 (
            .O(N__21850),
            .I(N__21837));
    Odrv4 I__3977 (
            .O(N__21847),
            .I(wrtrigmask_0));
    Odrv4 I__3976 (
            .O(N__21842),
            .I(wrtrigmask_0));
    Odrv4 I__3975 (
            .O(N__21837),
            .I(wrtrigmask_0));
    InMux I__3974 (
            .O(N__21830),
            .I(N__21826));
    InMux I__3973 (
            .O(N__21829),
            .I(N__21823));
    LocalMux I__3972 (
            .O(N__21826),
            .I(maskRegister_0));
    LocalMux I__3971 (
            .O(N__21823),
            .I(maskRegister_0));
    InMux I__3970 (
            .O(N__21818),
            .I(N__21811));
    InMux I__3969 (
            .O(N__21817),
            .I(N__21811));
    InMux I__3968 (
            .O(N__21816),
            .I(N__21808));
    LocalMux I__3967 (
            .O(N__21811),
            .I(N__21805));
    LocalMux I__3966 (
            .O(N__21808),
            .I(configRegister_20_adj_1382));
    Odrv4 I__3965 (
            .O(N__21805),
            .I(configRegister_20_adj_1382));
    InMux I__3964 (
            .O(N__21800),
            .I(N__21797));
    LocalMux I__3963 (
            .O(N__21797),
            .I(N__21793));
    InMux I__3962 (
            .O(N__21796),
            .I(N__21790));
    Odrv12 I__3961 (
            .O(N__21793),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6 ));
    LocalMux I__3960 (
            .O(N__21790),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6 ));
    CascadeMux I__3959 (
            .O(N__21785),
            .I(N__21782));
    InMux I__3958 (
            .O(N__21782),
            .I(N__21779));
    LocalMux I__3957 (
            .O(N__21779),
            .I(N__21776));
    Odrv4 I__3956 (
            .O(N__21776),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_7 ));
    CascadeMux I__3955 (
            .O(N__21773),
            .I(N__21770));
    InMux I__3954 (
            .O(N__21770),
            .I(N__21767));
    LocalMux I__3953 (
            .O(N__21767),
            .I(N__21763));
    InMux I__3952 (
            .O(N__21766),
            .I(N__21760));
    Odrv4 I__3951 (
            .O(N__21763),
            .I(configRegister_15_adj_1385));
    LocalMux I__3950 (
            .O(N__21760),
            .I(configRegister_15_adj_1385));
    InMux I__3949 (
            .O(N__21755),
            .I(N__21751));
    InMux I__3948 (
            .O(N__21754),
            .I(N__21748));
    LocalMux I__3947 (
            .O(N__21751),
            .I(configRegister_24_adj_1378));
    LocalMux I__3946 (
            .O(N__21748),
            .I(configRegister_24_adj_1378));
    CascadeMux I__3945 (
            .O(N__21743),
            .I(N__21738));
    CascadeMux I__3944 (
            .O(N__21742),
            .I(N__21735));
    InMux I__3943 (
            .O(N__21741),
            .I(N__21716));
    InMux I__3942 (
            .O(N__21738),
            .I(N__21716));
    InMux I__3941 (
            .O(N__21735),
            .I(N__21716));
    InMux I__3940 (
            .O(N__21734),
            .I(N__21716));
    InMux I__3939 (
            .O(N__21733),
            .I(N__21716));
    InMux I__3938 (
            .O(N__21732),
            .I(N__21716));
    InMux I__3937 (
            .O(N__21731),
            .I(N__21713));
    InMux I__3936 (
            .O(N__21730),
            .I(N__21708));
    InMux I__3935 (
            .O(N__21729),
            .I(N__21708));
    LocalMux I__3934 (
            .O(N__21716),
            .I(N__21705));
    LocalMux I__3933 (
            .O(N__21713),
            .I(N__21702));
    LocalMux I__3932 (
            .O(N__21708),
            .I(N__21699));
    Span4Mux_h I__3931 (
            .O(N__21705),
            .I(N__21694));
    Span4Mux_h I__3930 (
            .O(N__21702),
            .I(N__21694));
    Span4Mux_s3_h I__3929 (
            .O(N__21699),
            .I(N__21691));
    Span4Mux_v I__3928 (
            .O(N__21694),
            .I(N__21688));
    Odrv4 I__3927 (
            .O(N__21691),
            .I(\Inst_eia232.Inst_transmitter.n4246 ));
    Odrv4 I__3926 (
            .O(N__21688),
            .I(\Inst_eia232.Inst_transmitter.n4246 ));
    InMux I__3925 (
            .O(N__21683),
            .I(N__21678));
    CEMux I__3924 (
            .O(N__21682),
            .I(N__21673));
    InMux I__3923 (
            .O(N__21681),
            .I(N__21670));
    LocalMux I__3922 (
            .O(N__21678),
            .I(N__21659));
    CascadeMux I__3921 (
            .O(N__21677),
            .I(N__21652));
    CascadeMux I__3920 (
            .O(N__21676),
            .I(N__21649));
    LocalMux I__3919 (
            .O(N__21673),
            .I(N__21646));
    LocalMux I__3918 (
            .O(N__21670),
            .I(N__21643));
    InMux I__3917 (
            .O(N__21669),
            .I(N__21638));
    InMux I__3916 (
            .O(N__21668),
            .I(N__21638));
    InMux I__3915 (
            .O(N__21667),
            .I(N__21633));
    InMux I__3914 (
            .O(N__21666),
            .I(N__21633));
    InMux I__3913 (
            .O(N__21665),
            .I(N__21624));
    InMux I__3912 (
            .O(N__21664),
            .I(N__21624));
    InMux I__3911 (
            .O(N__21663),
            .I(N__21624));
    InMux I__3910 (
            .O(N__21662),
            .I(N__21624));
    Span4Mux_h I__3909 (
            .O(N__21659),
            .I(N__21621));
    CascadeMux I__3908 (
            .O(N__21658),
            .I(N__21618));
    CascadeMux I__3907 (
            .O(N__21657),
            .I(N__21615));
    CascadeMux I__3906 (
            .O(N__21656),
            .I(N__21612));
    CEMux I__3905 (
            .O(N__21655),
            .I(N__21607));
    InMux I__3904 (
            .O(N__21652),
            .I(N__21602));
    InMux I__3903 (
            .O(N__21649),
            .I(N__21602));
    Span4Mux_v I__3902 (
            .O(N__21646),
            .I(N__21599));
    Span4Mux_h I__3901 (
            .O(N__21643),
            .I(N__21596));
    LocalMux I__3900 (
            .O(N__21638),
            .I(N__21587));
    LocalMux I__3899 (
            .O(N__21633),
            .I(N__21587));
    LocalMux I__3898 (
            .O(N__21624),
            .I(N__21587));
    Span4Mux_v I__3897 (
            .O(N__21621),
            .I(N__21587));
    InMux I__3896 (
            .O(N__21618),
            .I(N__21584));
    InMux I__3895 (
            .O(N__21615),
            .I(N__21575));
    InMux I__3894 (
            .O(N__21612),
            .I(N__21575));
    InMux I__3893 (
            .O(N__21611),
            .I(N__21575));
    InMux I__3892 (
            .O(N__21610),
            .I(N__21575));
    LocalMux I__3891 (
            .O(N__21607),
            .I(N__21570));
    LocalMux I__3890 (
            .O(N__21602),
            .I(N__21570));
    Span4Mux_v I__3889 (
            .O(N__21599),
            .I(N__21565));
    Span4Mux_v I__3888 (
            .O(N__21596),
            .I(N__21565));
    Span4Mux_v I__3887 (
            .O(N__21587),
            .I(N__21562));
    LocalMux I__3886 (
            .O(N__21584),
            .I(n4005));
    LocalMux I__3885 (
            .O(N__21575),
            .I(n4005));
    Odrv12 I__3884 (
            .O(N__21570),
            .I(n4005));
    Odrv4 I__3883 (
            .O(N__21565),
            .I(n4005));
    Odrv4 I__3882 (
            .O(N__21562),
            .I(n4005));
    CascadeMux I__3881 (
            .O(N__21551),
            .I(N__21548));
    InMux I__3880 (
            .O(N__21548),
            .I(N__21542));
    InMux I__3879 (
            .O(N__21547),
            .I(N__21542));
    LocalMux I__3878 (
            .O(N__21542),
            .I(disabledGroupsReg_0));
    InMux I__3877 (
            .O(N__21539),
            .I(N__21536));
    LocalMux I__3876 (
            .O(N__21536),
            .I(N__21533));
    Span4Mux_s2_h I__3875 (
            .O(N__21533),
            .I(N__21529));
    InMux I__3874 (
            .O(N__21532),
            .I(N__21526));
    Span4Mux_h I__3873 (
            .O(N__21529),
            .I(N__21523));
    LocalMux I__3872 (
            .O(N__21526),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_0 ));
    Odrv4 I__3871 (
            .O(N__21523),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_0 ));
    InMux I__3870 (
            .O(N__21518),
            .I(N__21514));
    InMux I__3869 (
            .O(N__21517),
            .I(N__21511));
    LocalMux I__3868 (
            .O(N__21514),
            .I(configRegister_11_adj_1389));
    LocalMux I__3867 (
            .O(N__21511),
            .I(configRegister_11_adj_1389));
    InMux I__3866 (
            .O(N__21506),
            .I(N__21502));
    InMux I__3865 (
            .O(N__21505),
            .I(N__21499));
    LocalMux I__3864 (
            .O(N__21502),
            .I(configRegister_10_adj_1390));
    LocalMux I__3863 (
            .O(N__21499),
            .I(configRegister_10_adj_1390));
    CascadeMux I__3862 (
            .O(N__21494),
            .I(N__21491));
    InMux I__3861 (
            .O(N__21491),
            .I(N__21488));
    LocalMux I__3860 (
            .O(N__21488),
            .I(N__21484));
    InMux I__3859 (
            .O(N__21487),
            .I(N__21481));
    Span4Mux_v I__3858 (
            .O(N__21484),
            .I(N__21478));
    LocalMux I__3857 (
            .O(N__21481),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16 ));
    Odrv4 I__3856 (
            .O(N__21478),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16 ));
    InMux I__3855 (
            .O(N__21473),
            .I(N__21467));
    InMux I__3854 (
            .O(N__21472),
            .I(N__21467));
    LocalMux I__3853 (
            .O(N__21467),
            .I(N__21463));
    InMux I__3852 (
            .O(N__21466),
            .I(N__21460));
    Span4Mux_h I__3851 (
            .O(N__21463),
            .I(N__21457));
    LocalMux I__3850 (
            .O(N__21460),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16 ));
    Odrv4 I__3849 (
            .O(N__21457),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16 ));
    CascadeMux I__3848 (
            .O(N__21452),
            .I(N__21449));
    InMux I__3847 (
            .O(N__21449),
            .I(N__21445));
    InMux I__3846 (
            .O(N__21448),
            .I(N__21442));
    LocalMux I__3845 (
            .O(N__21445),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6 ));
    LocalMux I__3844 (
            .O(N__21442),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6 ));
    InMux I__3843 (
            .O(N__21437),
            .I(N__21433));
    InMux I__3842 (
            .O(N__21436),
            .I(N__21430));
    LocalMux I__3841 (
            .O(N__21433),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1 ));
    LocalMux I__3840 (
            .O(N__21430),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1 ));
    CascadeMux I__3839 (
            .O(N__21425),
            .I(N__21421));
    CascadeMux I__3838 (
            .O(N__21424),
            .I(N__21418));
    InMux I__3837 (
            .O(N__21421),
            .I(N__21415));
    InMux I__3836 (
            .O(N__21418),
            .I(N__21412));
    LocalMux I__3835 (
            .O(N__21415),
            .I(N__21409));
    LocalMux I__3834 (
            .O(N__21412),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4 ));
    Odrv4 I__3833 (
            .O(N__21409),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4 ));
    CascadeMux I__3832 (
            .O(N__21404),
            .I(N__21401));
    InMux I__3831 (
            .O(N__21401),
            .I(N__21397));
    InMux I__3830 (
            .O(N__21400),
            .I(N__21394));
    LocalMux I__3829 (
            .O(N__21397),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0 ));
    LocalMux I__3828 (
            .O(N__21394),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0 ));
    InMux I__3827 (
            .O(N__21389),
            .I(N__21386));
    LocalMux I__3826 (
            .O(N__21386),
            .I(N__21383));
    Span4Mux_h I__3825 (
            .O(N__21383),
            .I(N__21380));
    Odrv4 I__3824 (
            .O(N__21380),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n28 ));
    CascadeMux I__3823 (
            .O(N__21377),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n25_cascade_ ));
    InMux I__3822 (
            .O(N__21374),
            .I(N__21371));
    LocalMux I__3821 (
            .O(N__21371),
            .I(N__21368));
    Span4Mux_h I__3820 (
            .O(N__21368),
            .I(N__21365));
    Odrv4 I__3819 (
            .O(N__21365),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n27 ));
    CascadeMux I__3818 (
            .O(N__21362),
            .I(N__21359));
    InMux I__3817 (
            .O(N__21359),
            .I(N__21355));
    InMux I__3816 (
            .O(N__21358),
            .I(N__21352));
    LocalMux I__3815 (
            .O(N__21355),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13 ));
    LocalMux I__3814 (
            .O(N__21352),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13 ));
    InMux I__3813 (
            .O(N__21347),
            .I(N__21343));
    InMux I__3812 (
            .O(N__21346),
            .I(N__21340));
    LocalMux I__3811 (
            .O(N__21343),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3 ));
    LocalMux I__3810 (
            .O(N__21340),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3 ));
    CascadeMux I__3809 (
            .O(N__21335),
            .I(N__21331));
    InMux I__3808 (
            .O(N__21334),
            .I(N__21328));
    InMux I__3807 (
            .O(N__21331),
            .I(N__21325));
    LocalMux I__3806 (
            .O(N__21328),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5 ));
    LocalMux I__3805 (
            .O(N__21325),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5 ));
    InMux I__3804 (
            .O(N__21320),
            .I(N__21316));
    InMux I__3803 (
            .O(N__21319),
            .I(N__21313));
    LocalMux I__3802 (
            .O(N__21316),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8 ));
    LocalMux I__3801 (
            .O(N__21313),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8 ));
    InMux I__3800 (
            .O(N__21308),
            .I(N__21305));
    LocalMux I__3799 (
            .O(N__21305),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n26 ));
    InMux I__3798 (
            .O(N__21302),
            .I(N__21299));
    LocalMux I__3797 (
            .O(N__21299),
            .I(N__21295));
    InMux I__3796 (
            .O(N__21298),
            .I(N__21292));
    Odrv4 I__3795 (
            .O(N__21295),
            .I(valueRegister_6_adj_1370));
    LocalMux I__3794 (
            .O(N__21292),
            .I(valueRegister_6_adj_1370));
    InMux I__3793 (
            .O(N__21287),
            .I(N__21283));
    InMux I__3792 (
            .O(N__21286),
            .I(N__21280));
    LocalMux I__3791 (
            .O(N__21283),
            .I(configRegister_5_adj_1395));
    LocalMux I__3790 (
            .O(N__21280),
            .I(configRegister_5_adj_1395));
    InMux I__3789 (
            .O(N__21275),
            .I(N__21271));
    InMux I__3788 (
            .O(N__21274),
            .I(N__21268));
    LocalMux I__3787 (
            .O(N__21271),
            .I(valueRegister_7_adj_1369));
    LocalMux I__3786 (
            .O(N__21268),
            .I(valueRegister_7_adj_1369));
    InMux I__3785 (
            .O(N__21263),
            .I(N__21260));
    LocalMux I__3784 (
            .O(N__21260),
            .I(N__21256));
    InMux I__3783 (
            .O(N__21259),
            .I(N__21253));
    Span4Mux_h I__3782 (
            .O(N__21256),
            .I(N__21248));
    LocalMux I__3781 (
            .O(N__21253),
            .I(N__21248));
    Span4Mux_h I__3780 (
            .O(N__21248),
            .I(N__21245));
    Odrv4 I__3779 (
            .O(N__21245),
            .I(input_c_4));
    CascadeMux I__3778 (
            .O(N__21242),
            .I(N__21238));
    InMux I__3777 (
            .O(N__21241),
            .I(N__21235));
    InMux I__3776 (
            .O(N__21238),
            .I(N__21232));
    LocalMux I__3775 (
            .O(N__21235),
            .I(\Inst_core.Inst_sync.synchronizedInput180_4 ));
    LocalMux I__3774 (
            .O(N__21232),
            .I(\Inst_core.Inst_sync.synchronizedInput180_4 ));
    SRMux I__3773 (
            .O(N__21227),
            .I(N__21224));
    LocalMux I__3772 (
            .O(N__21224),
            .I(N__21221));
    Span4Mux_s2_v I__3771 (
            .O(N__21221),
            .I(N__21218));
    Odrv4 I__3770 (
            .O(N__21218),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4765 ));
    CascadeMux I__3769 (
            .O(N__21215),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n25_cascade_ ));
    InMux I__3768 (
            .O(N__21212),
            .I(N__21209));
    LocalMux I__3767 (
            .O(N__21209),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n27 ));
    InMux I__3766 (
            .O(N__21206),
            .I(N__21203));
    LocalMux I__3765 (
            .O(N__21203),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n26 ));
    SRMux I__3764 (
            .O(N__21200),
            .I(N__21197));
    LocalMux I__3763 (
            .O(N__21197),
            .I(N__21194));
    Span4Mux_v I__3762 (
            .O(N__21194),
            .I(N__21191));
    Span4Mux_h I__3761 (
            .O(N__21191),
            .I(N__21188));
    Odrv4 I__3760 (
            .O(N__21188),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4766 ));
    InMux I__3759 (
            .O(N__21185),
            .I(N__21182));
    LocalMux I__3758 (
            .O(N__21182),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n28 ));
    InMux I__3757 (
            .O(N__21179),
            .I(N__21175));
    InMux I__3756 (
            .O(N__21178),
            .I(N__21172));
    LocalMux I__3755 (
            .O(N__21175),
            .I(N__21169));
    LocalMux I__3754 (
            .O(N__21172),
            .I(\Inst_core.Inst_sync.filteredInput_5 ));
    Odrv4 I__3753 (
            .O(N__21169),
            .I(\Inst_core.Inst_sync.filteredInput_5 ));
    CascadeMux I__3752 (
            .O(N__21164),
            .I(\Inst_core.Inst_sync.n9063_cascade_ ));
    CascadeMux I__3751 (
            .O(N__21161),
            .I(N__21158));
    InMux I__3750 (
            .O(N__21158),
            .I(N__21155));
    LocalMux I__3749 (
            .O(N__21155),
            .I(syncedInput_5));
    InMux I__3748 (
            .O(N__21152),
            .I(N__21148));
    InMux I__3747 (
            .O(N__21151),
            .I(N__21145));
    LocalMux I__3746 (
            .O(N__21148),
            .I(N__21139));
    LocalMux I__3745 (
            .O(N__21145),
            .I(N__21139));
    InMux I__3744 (
            .O(N__21144),
            .I(N__21136));
    Odrv4 I__3743 (
            .O(N__21139),
            .I(\Inst_core.Inst_sync.synchronizedInput_4 ));
    LocalMux I__3742 (
            .O(N__21136),
            .I(\Inst_core.Inst_sync.synchronizedInput_4 ));
    InMux I__3741 (
            .O(N__21131),
            .I(N__21128));
    LocalMux I__3740 (
            .O(N__21128),
            .I(N__21125));
    Span4Mux_h I__3739 (
            .O(N__21125),
            .I(N__21121));
    InMux I__3738 (
            .O(N__21124),
            .I(N__21118));
    Span4Mux_s1_v I__3737 (
            .O(N__21121),
            .I(N__21115));
    LocalMux I__3736 (
            .O(N__21118),
            .I(\Inst_core.Inst_sync.filteredInput_4 ));
    Odrv4 I__3735 (
            .O(N__21115),
            .I(\Inst_core.Inst_sync.filteredInput_4 ));
    InMux I__3734 (
            .O(N__21110),
            .I(N__21106));
    InMux I__3733 (
            .O(N__21109),
            .I(N__21103));
    LocalMux I__3732 (
            .O(N__21106),
            .I(\Inst_core.Inst_sync.demuxedInput_4 ));
    LocalMux I__3731 (
            .O(N__21103),
            .I(\Inst_core.Inst_sync.demuxedInput_4 ));
    CascadeMux I__3730 (
            .O(N__21098),
            .I(\Inst_core.Inst_sync.n9057_cascade_ ));
    CascadeMux I__3729 (
            .O(N__21095),
            .I(N__21092));
    InMux I__3728 (
            .O(N__21092),
            .I(N__21089));
    LocalMux I__3727 (
            .O(N__21089),
            .I(syncedInput_4));
    InMux I__3726 (
            .O(N__21086),
            .I(N__21083));
    LocalMux I__3725 (
            .O(N__21083),
            .I(\Inst_core.Inst_sync.Inst_filter.input180Delay_6 ));
    SRMux I__3724 (
            .O(N__21080),
            .I(N__21077));
    LocalMux I__3723 (
            .O(N__21077),
            .I(N__21074));
    Span4Mux_h I__3722 (
            .O(N__21074),
            .I(N__21071));
    Span4Mux_v I__3721 (
            .O(N__21071),
            .I(N__21068));
    Odrv4 I__3720 (
            .O(N__21068),
            .I(\Inst_core.Inst_sync.Inst_filter.n4734 ));
    InMux I__3719 (
            .O(N__21065),
            .I(N__21062));
    LocalMux I__3718 (
            .O(N__21062),
            .I(\Inst_core.Inst_sync.Inst_filter.input180Delay_5 ));
    SRMux I__3717 (
            .O(N__21059),
            .I(N__21056));
    LocalMux I__3716 (
            .O(N__21056),
            .I(N__21053));
    Span4Mux_h I__3715 (
            .O(N__21053),
            .I(N__21050));
    Odrv4 I__3714 (
            .O(N__21050),
            .I(\Inst_core.Inst_sync.Inst_filter.n4733 ));
    CascadeMux I__3713 (
            .O(N__21047),
            .I(N__21044));
    InMux I__3712 (
            .O(N__21044),
            .I(N__21041));
    LocalMux I__3711 (
            .O(N__21041),
            .I(N__21037));
    InMux I__3710 (
            .O(N__21040),
            .I(N__21034));
    Span4Mux_v I__3709 (
            .O(N__21037),
            .I(N__21031));
    LocalMux I__3708 (
            .O(N__21034),
            .I(\Inst_core.Inst_sync.filteredInput_2 ));
    Odrv4 I__3707 (
            .O(N__21031),
            .I(\Inst_core.Inst_sync.filteredInput_2 ));
    CascadeMux I__3706 (
            .O(N__21026),
            .I(\Inst_core.Inst_sync.n2789_cascade_ ));
    CascadeMux I__3705 (
            .O(N__21023),
            .I(N__21020));
    InMux I__3704 (
            .O(N__21020),
            .I(N__21017));
    LocalMux I__3703 (
            .O(N__21017),
            .I(syncedInput_2));
    InMux I__3702 (
            .O(N__21014),
            .I(N__21011));
    LocalMux I__3701 (
            .O(N__21011),
            .I(N__21007));
    InMux I__3700 (
            .O(N__21010),
            .I(N__21004));
    Span4Mux_v I__3699 (
            .O(N__21007),
            .I(N__21001));
    LocalMux I__3698 (
            .O(N__21004),
            .I(\Inst_core.Inst_sync.demuxedInput_6 ));
    Odrv4 I__3697 (
            .O(N__21001),
            .I(\Inst_core.Inst_sync.demuxedInput_6 ));
    CascadeMux I__3696 (
            .O(N__20996),
            .I(N__20992));
    InMux I__3695 (
            .O(N__20995),
            .I(N__20989));
    InMux I__3694 (
            .O(N__20992),
            .I(N__20986));
    LocalMux I__3693 (
            .O(N__20989),
            .I(\Inst_core.Inst_sync.filteredInput_6 ));
    LocalMux I__3692 (
            .O(N__20986),
            .I(\Inst_core.Inst_sync.filteredInput_6 ));
    InMux I__3691 (
            .O(N__20981),
            .I(N__20977));
    InMux I__3690 (
            .O(N__20980),
            .I(N__20974));
    LocalMux I__3689 (
            .O(N__20977),
            .I(maskRegister_4_adj_1284));
    LocalMux I__3688 (
            .O(N__20974),
            .I(maskRegister_4_adj_1284));
    SRMux I__3687 (
            .O(N__20969),
            .I(N__20966));
    LocalMux I__3686 (
            .O(N__20966),
            .I(N__20963));
    Sp12to4 I__3685 (
            .O(N__20963),
            .I(N__20960));
    Odrv12 I__3684 (
            .O(N__20960),
            .I(\Inst_core.Inst_sync.Inst_filter.n4637 ));
    InMux I__3683 (
            .O(N__20957),
            .I(N__20953));
    InMux I__3682 (
            .O(N__20956),
            .I(N__20950));
    LocalMux I__3681 (
            .O(N__20953),
            .I(N__20947));
    LocalMux I__3680 (
            .O(N__20950),
            .I(maskRegister_1));
    Odrv12 I__3679 (
            .O(N__20947),
            .I(maskRegister_1));
    SRMux I__3678 (
            .O(N__20942),
            .I(N__20939));
    LocalMux I__3677 (
            .O(N__20939),
            .I(N__20936));
    Span4Mux_v I__3676 (
            .O(N__20936),
            .I(N__20933));
    Odrv4 I__3675 (
            .O(N__20933),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4739 ));
    InMux I__3674 (
            .O(N__20930),
            .I(N__20927));
    LocalMux I__3673 (
            .O(N__20927),
            .I(\Inst_core.Inst_sync.Inst_filter.input180Delay_7 ));
    InMux I__3672 (
            .O(N__20924),
            .I(N__20920));
    InMux I__3671 (
            .O(N__20923),
            .I(N__20917));
    LocalMux I__3670 (
            .O(N__20920),
            .I(N__20914));
    LocalMux I__3669 (
            .O(N__20917),
            .I(maskRegister_1_adj_1287));
    Odrv4 I__3668 (
            .O(N__20914),
            .I(maskRegister_1_adj_1287));
    InMux I__3667 (
            .O(N__20909),
            .I(N__20905));
    InMux I__3666 (
            .O(N__20908),
            .I(N__20902));
    LocalMux I__3665 (
            .O(N__20905),
            .I(maskRegister_2_adj_1286));
    LocalMux I__3664 (
            .O(N__20902),
            .I(maskRegister_2_adj_1286));
    InMux I__3663 (
            .O(N__20897),
            .I(N__20893));
    InMux I__3662 (
            .O(N__20896),
            .I(N__20890));
    LocalMux I__3661 (
            .O(N__20893),
            .I(N__20887));
    LocalMux I__3660 (
            .O(N__20890),
            .I(maskRegister_3_adj_1285));
    Odrv12 I__3659 (
            .O(N__20887),
            .I(maskRegister_3_adj_1285));
    InMux I__3658 (
            .O(N__20882),
            .I(N__20879));
    LocalMux I__3657 (
            .O(N__20879),
            .I(N__20875));
    InMux I__3656 (
            .O(N__20878),
            .I(N__20872));
    Span4Mux_v I__3655 (
            .O(N__20875),
            .I(N__20869));
    LocalMux I__3654 (
            .O(N__20872),
            .I(maskRegister_5_adj_1283));
    Odrv4 I__3653 (
            .O(N__20869),
            .I(maskRegister_5_adj_1283));
    InMux I__3652 (
            .O(N__20864),
            .I(N__20859));
    InMux I__3651 (
            .O(N__20863),
            .I(N__20854));
    InMux I__3650 (
            .O(N__20862),
            .I(N__20854));
    LocalMux I__3649 (
            .O(N__20859),
            .I(configRegister_20_adj_1302));
    LocalMux I__3648 (
            .O(N__20854),
            .I(configRegister_20_adj_1302));
    CascadeMux I__3647 (
            .O(N__20849),
            .I(N__20846));
    InMux I__3646 (
            .O(N__20846),
            .I(N__20842));
    InMux I__3645 (
            .O(N__20845),
            .I(N__20839));
    LocalMux I__3644 (
            .O(N__20842),
            .I(configRegister_24_adj_1298));
    LocalMux I__3643 (
            .O(N__20839),
            .I(configRegister_24_adj_1298));
    InMux I__3642 (
            .O(N__20834),
            .I(N__20830));
    InMux I__3641 (
            .O(N__20833),
            .I(N__20827));
    LocalMux I__3640 (
            .O(N__20830),
            .I(N__20824));
    LocalMux I__3639 (
            .O(N__20827),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16 ));
    Odrv4 I__3638 (
            .O(N__20824),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16 ));
    CascadeMux I__3637 (
            .O(N__20819),
            .I(N__20814));
    InMux I__3636 (
            .O(N__20818),
            .I(N__20809));
    InMux I__3635 (
            .O(N__20817),
            .I(N__20809));
    InMux I__3634 (
            .O(N__20814),
            .I(N__20806));
    LocalMux I__3633 (
            .O(N__20809),
            .I(N__20803));
    LocalMux I__3632 (
            .O(N__20806),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16 ));
    Odrv4 I__3631 (
            .O(N__20803),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16 ));
    InMux I__3630 (
            .O(N__20798),
            .I(N__20794));
    CascadeMux I__3629 (
            .O(N__20797),
            .I(N__20791));
    LocalMux I__3628 (
            .O(N__20794),
            .I(N__20787));
    InMux I__3627 (
            .O(N__20791),
            .I(N__20782));
    InMux I__3626 (
            .O(N__20790),
            .I(N__20782));
    Odrv12 I__3625 (
            .O(N__20787),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0 ));
    LocalMux I__3624 (
            .O(N__20782),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0 ));
    CascadeMux I__3623 (
            .O(N__20777),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_cascade_ ));
    InMux I__3622 (
            .O(N__20774),
            .I(N__20771));
    LocalMux I__3621 (
            .O(N__20771),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9078 ));
    CascadeMux I__3620 (
            .O(N__20768),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_cascade_ ));
    CascadeMux I__3619 (
            .O(N__20765),
            .I(N__20758));
    CascadeMux I__3618 (
            .O(N__20764),
            .I(N__20755));
    InMux I__3617 (
            .O(N__20763),
            .I(N__20752));
    InMux I__3616 (
            .O(N__20762),
            .I(N__20743));
    InMux I__3615 (
            .O(N__20761),
            .I(N__20743));
    InMux I__3614 (
            .O(N__20758),
            .I(N__20743));
    InMux I__3613 (
            .O(N__20755),
            .I(N__20743));
    LocalMux I__3612 (
            .O(N__20752),
            .I(configRegister_21_adj_1301));
    LocalMux I__3611 (
            .O(N__20743),
            .I(configRegister_21_adj_1301));
    InMux I__3610 (
            .O(N__20738),
            .I(N__20733));
    InMux I__3609 (
            .O(N__20737),
            .I(N__20728));
    InMux I__3608 (
            .O(N__20736),
            .I(N__20728));
    LocalMux I__3607 (
            .O(N__20733),
            .I(configRegister_23_adj_1299));
    LocalMux I__3606 (
            .O(N__20728),
            .I(configRegister_23_adj_1299));
    InMux I__3605 (
            .O(N__20723),
            .I(N__20716));
    InMux I__3604 (
            .O(N__20722),
            .I(N__20716));
    InMux I__3603 (
            .O(N__20721),
            .I(N__20713));
    LocalMux I__3602 (
            .O(N__20716),
            .I(N__20710));
    LocalMux I__3601 (
            .O(N__20713),
            .I(configRegister_22_adj_1300));
    Odrv4 I__3600 (
            .O(N__20710),
            .I(configRegister_22_adj_1300));
    CascadeMux I__3599 (
            .O(N__20705),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9072_cascade_ ));
    InMux I__3598 (
            .O(N__20702),
            .I(N__20696));
    InMux I__3597 (
            .O(N__20701),
            .I(N__20692));
    InMux I__3596 (
            .O(N__20700),
            .I(N__20684));
    InMux I__3595 (
            .O(N__20699),
            .I(N__20684));
    LocalMux I__3594 (
            .O(N__20696),
            .I(N__20681));
    InMux I__3593 (
            .O(N__20695),
            .I(N__20678));
    LocalMux I__3592 (
            .O(N__20692),
            .I(N__20675));
    InMux I__3591 (
            .O(N__20691),
            .I(N__20672));
    CascadeMux I__3590 (
            .O(N__20690),
            .I(N__20669));
    InMux I__3589 (
            .O(N__20689),
            .I(N__20666));
    LocalMux I__3588 (
            .O(N__20684),
            .I(N__20663));
    Span4Mux_v I__3587 (
            .O(N__20681),
            .I(N__20654));
    LocalMux I__3586 (
            .O(N__20678),
            .I(N__20654));
    Span4Mux_s3_v I__3585 (
            .O(N__20675),
            .I(N__20654));
    LocalMux I__3584 (
            .O(N__20672),
            .I(N__20654));
    InMux I__3583 (
            .O(N__20669),
            .I(N__20651));
    LocalMux I__3582 (
            .O(N__20666),
            .I(N__20644));
    Span4Mux_v I__3581 (
            .O(N__20663),
            .I(N__20644));
    Span4Mux_v I__3580 (
            .O(N__20654),
            .I(N__20644));
    LocalMux I__3579 (
            .O(N__20651),
            .I(N__20641));
    Span4Mux_v I__3578 (
            .O(N__20644),
            .I(N__20638));
    Odrv4 I__3577 (
            .O(N__20641),
            .I(wrtrigval_0));
    Odrv4 I__3576 (
            .O(N__20638),
            .I(wrtrigval_0));
    InMux I__3575 (
            .O(N__20633),
            .I(N__20630));
    LocalMux I__3574 (
            .O(N__20630),
            .I(N__20625));
    InMux I__3573 (
            .O(N__20629),
            .I(N__20620));
    InMux I__3572 (
            .O(N__20628),
            .I(N__20620));
    Odrv4 I__3571 (
            .O(N__20625),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1 ));
    LocalMux I__3570 (
            .O(N__20620),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1 ));
    InMux I__3569 (
            .O(N__20615),
            .I(N__20611));
    InMux I__3568 (
            .O(N__20614),
            .I(N__20608));
    LocalMux I__3567 (
            .O(N__20611),
            .I(valueRegister_1));
    LocalMux I__3566 (
            .O(N__20608),
            .I(valueRegister_1));
    InMux I__3565 (
            .O(N__20603),
            .I(N__20599));
    CascadeMux I__3564 (
            .O(N__20602),
            .I(N__20594));
    LocalMux I__3563 (
            .O(N__20599),
            .I(N__20590));
    InMux I__3562 (
            .O(N__20598),
            .I(N__20587));
    InMux I__3561 (
            .O(N__20597),
            .I(N__20584));
    InMux I__3560 (
            .O(N__20594),
            .I(N__20581));
    CascadeMux I__3559 (
            .O(N__20593),
            .I(N__20577));
    Span4Mux_s2_v I__3558 (
            .O(N__20590),
            .I(N__20571));
    LocalMux I__3557 (
            .O(N__20587),
            .I(N__20571));
    LocalMux I__3556 (
            .O(N__20584),
            .I(N__20568));
    LocalMux I__3555 (
            .O(N__20581),
            .I(N__20565));
    InMux I__3554 (
            .O(N__20580),
            .I(N__20562));
    InMux I__3553 (
            .O(N__20577),
            .I(N__20558));
    InMux I__3552 (
            .O(N__20576),
            .I(N__20555));
    Span4Mux_v I__3551 (
            .O(N__20571),
            .I(N__20551));
    Span4Mux_v I__3550 (
            .O(N__20568),
            .I(N__20546));
    Span4Mux_v I__3549 (
            .O(N__20565),
            .I(N__20546));
    LocalMux I__3548 (
            .O(N__20562),
            .I(N__20543));
    InMux I__3547 (
            .O(N__20561),
            .I(N__20540));
    LocalMux I__3546 (
            .O(N__20558),
            .I(N__20535));
    LocalMux I__3545 (
            .O(N__20555),
            .I(N__20535));
    InMux I__3544 (
            .O(N__20554),
            .I(N__20532));
    Odrv4 I__3543 (
            .O(N__20551),
            .I(configRegister_26));
    Odrv4 I__3542 (
            .O(N__20546),
            .I(configRegister_26));
    Odrv12 I__3541 (
            .O(N__20543),
            .I(configRegister_26));
    LocalMux I__3540 (
            .O(N__20540),
            .I(configRegister_26));
    Odrv4 I__3539 (
            .O(N__20535),
            .I(configRegister_26));
    LocalMux I__3538 (
            .O(N__20532),
            .I(configRegister_26));
    InMux I__3537 (
            .O(N__20519),
            .I(N__20516));
    LocalMux I__3536 (
            .O(N__20516),
            .I(N__20513));
    Span4Mux_v I__3535 (
            .O(N__20513),
            .I(N__20510));
    Odrv4 I__3534 (
            .O(N__20510),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_1 ));
    InMux I__3533 (
            .O(N__20507),
            .I(N__20504));
    LocalMux I__3532 (
            .O(N__20504),
            .I(N__20501));
    Odrv4 I__3531 (
            .O(N__20501),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_3 ));
    InMux I__3530 (
            .O(N__20498),
            .I(N__20494));
    InMux I__3529 (
            .O(N__20497),
            .I(N__20491));
    LocalMux I__3528 (
            .O(N__20494),
            .I(N__20488));
    LocalMux I__3527 (
            .O(N__20491),
            .I(configRegister_0_adj_1400));
    Odrv12 I__3526 (
            .O(N__20488),
            .I(configRegister_0_adj_1400));
    InMux I__3525 (
            .O(N__20483),
            .I(N__20476));
    InMux I__3524 (
            .O(N__20482),
            .I(N__20476));
    InMux I__3523 (
            .O(N__20481),
            .I(N__20473));
    LocalMux I__3522 (
            .O(N__20476),
            .I(N__20470));
    LocalMux I__3521 (
            .O(N__20473),
            .I(configRegister_20_adj_1342));
    Odrv4 I__3520 (
            .O(N__20470),
            .I(configRegister_20_adj_1342));
    InMux I__3519 (
            .O(N__20465),
            .I(N__20462));
    LocalMux I__3518 (
            .O(N__20462),
            .I(N__20458));
    InMux I__3517 (
            .O(N__20461),
            .I(N__20455));
    Span4Mux_s3_v I__3516 (
            .O(N__20458),
            .I(N__20452));
    LocalMux I__3515 (
            .O(N__20455),
            .I(configRegister_4_adj_1396));
    Odrv4 I__3514 (
            .O(N__20452),
            .I(configRegister_4_adj_1396));
    CascadeMux I__3513 (
            .O(N__20447),
            .I(N__20442));
    InMux I__3512 (
            .O(N__20446),
            .I(N__20439));
    InMux I__3511 (
            .O(N__20445),
            .I(N__20436));
    InMux I__3510 (
            .O(N__20442),
            .I(N__20433));
    LocalMux I__3509 (
            .O(N__20439),
            .I(N__20428));
    LocalMux I__3508 (
            .O(N__20436),
            .I(N__20428));
    LocalMux I__3507 (
            .O(N__20433),
            .I(cmd_39));
    Odrv4 I__3506 (
            .O(N__20428),
            .I(cmd_39));
    SRMux I__3505 (
            .O(N__20423),
            .I(N__20420));
    LocalMux I__3504 (
            .O(N__20420),
            .I(N__20417));
    Odrv12 I__3503 (
            .O(N__20417),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4641 ));
    CascadeMux I__3502 (
            .O(N__20414),
            .I(N__20407));
    InMux I__3501 (
            .O(N__20413),
            .I(N__20404));
    InMux I__3500 (
            .O(N__20412),
            .I(N__20395));
    InMux I__3499 (
            .O(N__20411),
            .I(N__20395));
    InMux I__3498 (
            .O(N__20410),
            .I(N__20395));
    InMux I__3497 (
            .O(N__20407),
            .I(N__20395));
    LocalMux I__3496 (
            .O(N__20404),
            .I(configRegister_21_adj_1381));
    LocalMux I__3495 (
            .O(N__20395),
            .I(configRegister_21_adj_1381));
    InMux I__3494 (
            .O(N__20390),
            .I(N__20386));
    InMux I__3493 (
            .O(N__20389),
            .I(N__20383));
    LocalMux I__3492 (
            .O(N__20386),
            .I(maskRegister_6_adj_1362));
    LocalMux I__3491 (
            .O(N__20383),
            .I(maskRegister_6_adj_1362));
    InMux I__3490 (
            .O(N__20378),
            .I(N__20374));
    InMux I__3489 (
            .O(N__20377),
            .I(N__20371));
    LocalMux I__3488 (
            .O(N__20374),
            .I(maskRegister_7_adj_1361));
    LocalMux I__3487 (
            .O(N__20371),
            .I(maskRegister_7_adj_1361));
    InMux I__3486 (
            .O(N__20366),
            .I(N__20362));
    InMux I__3485 (
            .O(N__20365),
            .I(N__20359));
    LocalMux I__3484 (
            .O(N__20362),
            .I(maskRegister_4_adj_1364));
    LocalMux I__3483 (
            .O(N__20359),
            .I(maskRegister_4_adj_1364));
    InMux I__3482 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__3481 (
            .O(N__20351),
            .I(N__20348));
    Span4Mux_s2_v I__3480 (
            .O(N__20348),
            .I(N__20344));
    InMux I__3479 (
            .O(N__20347),
            .I(N__20341));
    Odrv4 I__3478 (
            .O(N__20344),
            .I(configRegister_6_adj_1394));
    LocalMux I__3477 (
            .O(N__20341),
            .I(configRegister_6_adj_1394));
    InMux I__3476 (
            .O(N__20336),
            .I(N__20332));
    InMux I__3475 (
            .O(N__20335),
            .I(N__20329));
    LocalMux I__3474 (
            .O(N__20332),
            .I(maskRegister_3_adj_1365));
    LocalMux I__3473 (
            .O(N__20329),
            .I(maskRegister_3_adj_1365));
    InMux I__3472 (
            .O(N__20324),
            .I(N__20321));
    LocalMux I__3471 (
            .O(N__20321),
            .I(N__20317));
    InMux I__3470 (
            .O(N__20320),
            .I(N__20314));
    Odrv4 I__3469 (
            .O(N__20317),
            .I(configRegister_7_adj_1393));
    LocalMux I__3468 (
            .O(N__20314),
            .I(configRegister_7_adj_1393));
    InMux I__3467 (
            .O(N__20309),
            .I(N__20306));
    LocalMux I__3466 (
            .O(N__20306),
            .I(N__20303));
    Span4Mux_s3_h I__3465 (
            .O(N__20303),
            .I(N__20300));
    Span4Mux_v I__3464 (
            .O(N__20300),
            .I(N__20296));
    InMux I__3463 (
            .O(N__20299),
            .I(N__20293));
    Odrv4 I__3462 (
            .O(N__20296),
            .I(valueRegister_0_adj_1296));
    LocalMux I__3461 (
            .O(N__20293),
            .I(valueRegister_0_adj_1296));
    CascadeMux I__3460 (
            .O(N__20288),
            .I(N__20285));
    InMux I__3459 (
            .O(N__20285),
            .I(N__20281));
    InMux I__3458 (
            .O(N__20284),
            .I(N__20278));
    LocalMux I__3457 (
            .O(N__20281),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11 ));
    LocalMux I__3456 (
            .O(N__20278),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11 ));
    InMux I__3455 (
            .O(N__20273),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7924 ));
    InMux I__3454 (
            .O(N__20270),
            .I(N__20266));
    InMux I__3453 (
            .O(N__20269),
            .I(N__20263));
    LocalMux I__3452 (
            .O(N__20266),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12 ));
    LocalMux I__3451 (
            .O(N__20263),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12 ));
    InMux I__3450 (
            .O(N__20258),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7925 ));
    InMux I__3449 (
            .O(N__20255),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7926 ));
    InMux I__3448 (
            .O(N__20252),
            .I(N__20248));
    InMux I__3447 (
            .O(N__20251),
            .I(N__20245));
    LocalMux I__3446 (
            .O(N__20248),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14 ));
    LocalMux I__3445 (
            .O(N__20245),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14 ));
    InMux I__3444 (
            .O(N__20240),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7927 ));
    InMux I__3443 (
            .O(N__20237),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7928 ));
    CascadeMux I__3442 (
            .O(N__20234),
            .I(N__20230));
    InMux I__3441 (
            .O(N__20233),
            .I(N__20227));
    InMux I__3440 (
            .O(N__20230),
            .I(N__20224));
    LocalMux I__3439 (
            .O(N__20227),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15 ));
    LocalMux I__3438 (
            .O(N__20224),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15 ));
    InMux I__3437 (
            .O(N__20219),
            .I(N__20216));
    LocalMux I__3436 (
            .O(N__20216),
            .I(N__20213));
    Span4Mux_v I__3435 (
            .O(N__20213),
            .I(N__20206));
    InMux I__3434 (
            .O(N__20212),
            .I(N__20201));
    InMux I__3433 (
            .O(N__20211),
            .I(N__20201));
    InMux I__3432 (
            .O(N__20210),
            .I(N__20198));
    InMux I__3431 (
            .O(N__20209),
            .I(N__20195));
    Odrv4 I__3430 (
            .O(N__20206),
            .I(\Inst_eia232.Inst_receiver.n7_adj_1264 ));
    LocalMux I__3429 (
            .O(N__20201),
            .I(\Inst_eia232.Inst_receiver.n7_adj_1264 ));
    LocalMux I__3428 (
            .O(N__20198),
            .I(\Inst_eia232.Inst_receiver.n7_adj_1264 ));
    LocalMux I__3427 (
            .O(N__20195),
            .I(\Inst_eia232.Inst_receiver.n7_adj_1264 ));
    InMux I__3426 (
            .O(N__20186),
            .I(N__20178));
    InMux I__3425 (
            .O(N__20185),
            .I(N__20165));
    InMux I__3424 (
            .O(N__20184),
            .I(N__20165));
    InMux I__3423 (
            .O(N__20183),
            .I(N__20165));
    InMux I__3422 (
            .O(N__20182),
            .I(N__20165));
    InMux I__3421 (
            .O(N__20181),
            .I(N__20165));
    LocalMux I__3420 (
            .O(N__20178),
            .I(N__20159));
    InMux I__3419 (
            .O(N__20177),
            .I(N__20154));
    InMux I__3418 (
            .O(N__20176),
            .I(N__20154));
    LocalMux I__3417 (
            .O(N__20165),
            .I(N__20151));
    InMux I__3416 (
            .O(N__20164),
            .I(N__20144));
    InMux I__3415 (
            .O(N__20163),
            .I(N__20144));
    InMux I__3414 (
            .O(N__20162),
            .I(N__20144));
    Odrv4 I__3413 (
            .O(N__20159),
            .I(\Inst_eia232.Inst_receiver.n957 ));
    LocalMux I__3412 (
            .O(N__20154),
            .I(\Inst_eia232.Inst_receiver.n957 ));
    Odrv4 I__3411 (
            .O(N__20151),
            .I(\Inst_eia232.Inst_receiver.n957 ));
    LocalMux I__3410 (
            .O(N__20144),
            .I(\Inst_eia232.Inst_receiver.n957 ));
    CascadeMux I__3409 (
            .O(N__20135),
            .I(N__20130));
    InMux I__3408 (
            .O(N__20134),
            .I(N__20123));
    InMux I__3407 (
            .O(N__20133),
            .I(N__20123));
    InMux I__3406 (
            .O(N__20130),
            .I(N__20116));
    InMux I__3405 (
            .O(N__20129),
            .I(N__20116));
    InMux I__3404 (
            .O(N__20128),
            .I(N__20116));
    LocalMux I__3403 (
            .O(N__20123),
            .I(N__20110));
    LocalMux I__3402 (
            .O(N__20116),
            .I(N__20110));
    InMux I__3401 (
            .O(N__20115),
            .I(N__20107));
    Span4Mux_h I__3400 (
            .O(N__20110),
            .I(N__20104));
    LocalMux I__3399 (
            .O(N__20107),
            .I(\Inst_eia232.Inst_receiver.bytecount_0 ));
    Odrv4 I__3398 (
            .O(N__20104),
            .I(\Inst_eia232.Inst_receiver.bytecount_0 ));
    CEMux I__3397 (
            .O(N__20099),
            .I(N__20095));
    CEMux I__3396 (
            .O(N__20098),
            .I(N__20092));
    LocalMux I__3395 (
            .O(N__20095),
            .I(N__20088));
    LocalMux I__3394 (
            .O(N__20092),
            .I(N__20085));
    InMux I__3393 (
            .O(N__20091),
            .I(N__20082));
    Span4Mux_h I__3392 (
            .O(N__20088),
            .I(N__20079));
    Span4Mux_s1_v I__3391 (
            .O(N__20085),
            .I(N__20076));
    LocalMux I__3390 (
            .O(N__20082),
            .I(N__20073));
    Span4Mux_v I__3389 (
            .O(N__20079),
            .I(N__20070));
    Span4Mux_v I__3388 (
            .O(N__20076),
            .I(N__20065));
    Span4Mux_h I__3387 (
            .O(N__20073),
            .I(N__20065));
    Odrv4 I__3386 (
            .O(N__20070),
            .I(\Inst_eia232.Inst_receiver.n3557 ));
    Odrv4 I__3385 (
            .O(N__20065),
            .I(\Inst_eia232.Inst_receiver.n3557 ));
    SRMux I__3384 (
            .O(N__20060),
            .I(N__20057));
    LocalMux I__3383 (
            .O(N__20057),
            .I(\Inst_eia232.Inst_receiver.n8376 ));
    InMux I__3382 (
            .O(N__20054),
            .I(N__20050));
    InMux I__3381 (
            .O(N__20053),
            .I(N__20047));
    LocalMux I__3380 (
            .O(N__20050),
            .I(configRegister_3_adj_1397));
    LocalMux I__3379 (
            .O(N__20047),
            .I(configRegister_3_adj_1397));
    InMux I__3378 (
            .O(N__20042),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7916 ));
    InMux I__3377 (
            .O(N__20039),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7917 ));
    InMux I__3376 (
            .O(N__20036),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7918 ));
    InMux I__3375 (
            .O(N__20033),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7919 ));
    CascadeMux I__3374 (
            .O(N__20030),
            .I(N__20026));
    InMux I__3373 (
            .O(N__20029),
            .I(N__20023));
    InMux I__3372 (
            .O(N__20026),
            .I(N__20020));
    LocalMux I__3371 (
            .O(N__20023),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7 ));
    LocalMux I__3370 (
            .O(N__20020),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7 ));
    InMux I__3369 (
            .O(N__20015),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7920 ));
    InMux I__3368 (
            .O(N__20012),
            .I(N__20008));
    InMux I__3367 (
            .O(N__20011),
            .I(N__20005));
    LocalMux I__3366 (
            .O(N__20008),
            .I(N__20002));
    LocalMux I__3365 (
            .O(N__20005),
            .I(configRegister_8_adj_1392));
    Odrv12 I__3364 (
            .O(N__20002),
            .I(configRegister_8_adj_1392));
    InMux I__3363 (
            .O(N__19997),
            .I(bfn_6_4_0_));
    CascadeMux I__3362 (
            .O(N__19994),
            .I(N__19991));
    InMux I__3361 (
            .O(N__19991),
            .I(N__19987));
    InMux I__3360 (
            .O(N__19990),
            .I(N__19984));
    LocalMux I__3359 (
            .O(N__19987),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9 ));
    LocalMux I__3358 (
            .O(N__19984),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9 ));
    InMux I__3357 (
            .O(N__19979),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7922 ));
    InMux I__3356 (
            .O(N__19976),
            .I(N__19972));
    InMux I__3355 (
            .O(N__19975),
            .I(N__19969));
    LocalMux I__3354 (
            .O(N__19972),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10 ));
    LocalMux I__3353 (
            .O(N__19969),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10 ));
    InMux I__3352 (
            .O(N__19964),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7923 ));
    InMux I__3351 (
            .O(N__19961),
            .I(bfn_6_3_0_));
    InMux I__3350 (
            .O(N__19958),
            .I(N__19954));
    InMux I__3349 (
            .O(N__19957),
            .I(N__19951));
    LocalMux I__3348 (
            .O(N__19954),
            .I(configRegister_1_adj_1399));
    LocalMux I__3347 (
            .O(N__19951),
            .I(configRegister_1_adj_1399));
    InMux I__3346 (
            .O(N__19946),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7914 ));
    InMux I__3345 (
            .O(N__19943),
            .I(N__19940));
    LocalMux I__3344 (
            .O(N__19940),
            .I(N__19936));
    InMux I__3343 (
            .O(N__19939),
            .I(N__19933));
    Odrv4 I__3342 (
            .O(N__19936),
            .I(configRegister_2_adj_1398));
    LocalMux I__3341 (
            .O(N__19933),
            .I(configRegister_2_adj_1398));
    CascadeMux I__3340 (
            .O(N__19928),
            .I(N__19925));
    InMux I__3339 (
            .O(N__19925),
            .I(N__19921));
    InMux I__3338 (
            .O(N__19924),
            .I(N__19918));
    LocalMux I__3337 (
            .O(N__19921),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2 ));
    LocalMux I__3336 (
            .O(N__19918),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2 ));
    InMux I__3335 (
            .O(N__19913),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7915 ));
    IoInMux I__3334 (
            .O(N__19910),
            .I(N__19907));
    LocalMux I__3333 (
            .O(N__19907),
            .I(N__19904));
    Span4Mux_s0_v I__3332 (
            .O(N__19904),
            .I(N__19900));
    InMux I__3331 (
            .O(N__19903),
            .I(N__19897));
    Odrv4 I__3330 (
            .O(N__19900),
            .I(testcnt_c_1));
    LocalMux I__3329 (
            .O(N__19897),
            .I(testcnt_c_1));
    InMux I__3328 (
            .O(N__19892),
            .I(n7862));
    IoInMux I__3327 (
            .O(N__19889),
            .I(N__19886));
    LocalMux I__3326 (
            .O(N__19886),
            .I(N__19883));
    IoSpan4Mux I__3325 (
            .O(N__19883),
            .I(N__19879));
    InMux I__3324 (
            .O(N__19882),
            .I(N__19876));
    Odrv4 I__3323 (
            .O(N__19879),
            .I(testcnt_c_2));
    LocalMux I__3322 (
            .O(N__19876),
            .I(testcnt_c_2));
    InMux I__3321 (
            .O(N__19871),
            .I(n7863));
    IoInMux I__3320 (
            .O(N__19868),
            .I(N__19864));
    InMux I__3319 (
            .O(N__19867),
            .I(N__19861));
    LocalMux I__3318 (
            .O(N__19864),
            .I(testcnt_c_3));
    LocalMux I__3317 (
            .O(N__19861),
            .I(testcnt_c_3));
    InMux I__3316 (
            .O(N__19856),
            .I(n7864));
    IoInMux I__3315 (
            .O(N__19853),
            .I(N__19849));
    InMux I__3314 (
            .O(N__19852),
            .I(N__19846));
    LocalMux I__3313 (
            .O(N__19849),
            .I(testcnt_c_4));
    LocalMux I__3312 (
            .O(N__19846),
            .I(testcnt_c_4));
    InMux I__3311 (
            .O(N__19841),
            .I(n7865));
    IoInMux I__3310 (
            .O(N__19838),
            .I(N__19834));
    InMux I__3309 (
            .O(N__19837),
            .I(N__19831));
    LocalMux I__3308 (
            .O(N__19834),
            .I(testcnt_c_5));
    LocalMux I__3307 (
            .O(N__19831),
            .I(testcnt_c_5));
    InMux I__3306 (
            .O(N__19826),
            .I(n7866));
    IoInMux I__3305 (
            .O(N__19823),
            .I(N__19820));
    LocalMux I__3304 (
            .O(N__19820),
            .I(N__19817));
    Span4Mux_s0_v I__3303 (
            .O(N__19817),
            .I(N__19813));
    InMux I__3302 (
            .O(N__19816),
            .I(N__19810));
    Odrv4 I__3301 (
            .O(N__19813),
            .I(testcnt_c_6));
    LocalMux I__3300 (
            .O(N__19810),
            .I(testcnt_c_6));
    InMux I__3299 (
            .O(N__19805),
            .I(n7867));
    InMux I__3298 (
            .O(N__19802),
            .I(n7868));
    IoInMux I__3297 (
            .O(N__19799),
            .I(N__19796));
    LocalMux I__3296 (
            .O(N__19796),
            .I(N__19793));
    Span4Mux_s0_v I__3295 (
            .O(N__19793),
            .I(N__19789));
    InMux I__3294 (
            .O(N__19792),
            .I(N__19786));
    Odrv4 I__3293 (
            .O(N__19789),
            .I(testcnt_c_7));
    LocalMux I__3292 (
            .O(N__19786),
            .I(testcnt_c_7));
    InMux I__3291 (
            .O(N__19781),
            .I(N__19778));
    LocalMux I__3290 (
            .O(N__19778),
            .I(N__19775));
    Span4Mux_s2_v I__3289 (
            .O(N__19775),
            .I(N__19771));
    InMux I__3288 (
            .O(N__19774),
            .I(N__19768));
    Span4Mux_v I__3287 (
            .O(N__19771),
            .I(N__19763));
    LocalMux I__3286 (
            .O(N__19768),
            .I(N__19763));
    Span4Mux_h I__3285 (
            .O(N__19763),
            .I(N__19760));
    Odrv4 I__3284 (
            .O(N__19760),
            .I(\GENERIC_FIFO_1.n8819 ));
    InMux I__3283 (
            .O(N__19757),
            .I(N__19753));
    InMux I__3282 (
            .O(N__19756),
            .I(N__19749));
    LocalMux I__3281 (
            .O(N__19753),
            .I(N__19746));
    InMux I__3280 (
            .O(N__19752),
            .I(N__19742));
    LocalMux I__3279 (
            .O(N__19749),
            .I(N__19736));
    Span4Mux_h I__3278 (
            .O(N__19746),
            .I(N__19736));
    InMux I__3277 (
            .O(N__19745),
            .I(N__19733));
    LocalMux I__3276 (
            .O(N__19742),
            .I(N__19730));
    InMux I__3275 (
            .O(N__19741),
            .I(N__19726));
    Span4Mux_v I__3274 (
            .O(N__19736),
            .I(N__19721));
    LocalMux I__3273 (
            .O(N__19733),
            .I(N__19721));
    Span4Mux_h I__3272 (
            .O(N__19730),
            .I(N__19718));
    InMux I__3271 (
            .O(N__19729),
            .I(N__19715));
    LocalMux I__3270 (
            .O(N__19726),
            .I(\GENERIC_FIFO_1.read_pointer_7 ));
    Odrv4 I__3269 (
            .O(N__19721),
            .I(\GENERIC_FIFO_1.read_pointer_7 ));
    Odrv4 I__3268 (
            .O(N__19718),
            .I(\GENERIC_FIFO_1.read_pointer_7 ));
    LocalMux I__3267 (
            .O(N__19715),
            .I(\GENERIC_FIFO_1.read_pointer_7 ));
    InMux I__3266 (
            .O(N__19706),
            .I(N__19701));
    InMux I__3265 (
            .O(N__19705),
            .I(N__19695));
    InMux I__3264 (
            .O(N__19704),
            .I(N__19695));
    LocalMux I__3263 (
            .O(N__19701),
            .I(N__19692));
    InMux I__3262 (
            .O(N__19700),
            .I(N__19679));
    LocalMux I__3261 (
            .O(N__19695),
            .I(N__19676));
    Span4Mux_h I__3260 (
            .O(N__19692),
            .I(N__19673));
    InMux I__3259 (
            .O(N__19691),
            .I(N__19668));
    InMux I__3258 (
            .O(N__19690),
            .I(N__19668));
    InMux I__3257 (
            .O(N__19689),
            .I(N__19649));
    InMux I__3256 (
            .O(N__19688),
            .I(N__19649));
    InMux I__3255 (
            .O(N__19687),
            .I(N__19649));
    InMux I__3254 (
            .O(N__19686),
            .I(N__19649));
    InMux I__3253 (
            .O(N__19685),
            .I(N__19649));
    InMux I__3252 (
            .O(N__19684),
            .I(N__19649));
    InMux I__3251 (
            .O(N__19683),
            .I(N__19649));
    InMux I__3250 (
            .O(N__19682),
            .I(N__19646));
    LocalMux I__3249 (
            .O(N__19679),
            .I(N__19641));
    Span4Mux_v I__3248 (
            .O(N__19676),
            .I(N__19641));
    Span4Mux_v I__3247 (
            .O(N__19673),
            .I(N__19636));
    LocalMux I__3246 (
            .O(N__19668),
            .I(N__19636));
    InMux I__3245 (
            .O(N__19667),
            .I(N__19627));
    InMux I__3244 (
            .O(N__19666),
            .I(N__19627));
    InMux I__3243 (
            .O(N__19665),
            .I(N__19627));
    InMux I__3242 (
            .O(N__19664),
            .I(N__19627));
    LocalMux I__3241 (
            .O(N__19649),
            .I(N__19624));
    LocalMux I__3240 (
            .O(N__19646),
            .I(N__19619));
    IoSpan4Mux I__3239 (
            .O(N__19641),
            .I(N__19619));
    Span4Mux_h I__3238 (
            .O(N__19636),
            .I(N__19616));
    LocalMux I__3237 (
            .O(N__19627),
            .I(N__19613));
    Span4Mux_h I__3236 (
            .O(N__19624),
            .I(N__19605));
    Span4Mux_s1_v I__3235 (
            .O(N__19619),
            .I(N__19605));
    Span4Mux_v I__3234 (
            .O(N__19616),
            .I(N__19605));
    Span4Mux_h I__3233 (
            .O(N__19613),
            .I(N__19602));
    InMux I__3232 (
            .O(N__19612),
            .I(N__19599));
    Odrv4 I__3231 (
            .O(N__19605),
            .I(\GENERIC_FIFO_1.n141 ));
    Odrv4 I__3230 (
            .O(N__19602),
            .I(\GENERIC_FIFO_1.n141 ));
    LocalMux I__3229 (
            .O(N__19599),
            .I(\GENERIC_FIFO_1.n141 ));
    InMux I__3228 (
            .O(N__19592),
            .I(N__19589));
    LocalMux I__3227 (
            .O(N__19589),
            .I(N__19585));
    InMux I__3226 (
            .O(N__19588),
            .I(N__19582));
    Span4Mux_v I__3225 (
            .O(N__19585),
            .I(N__19579));
    LocalMux I__3224 (
            .O(N__19582),
            .I(N__19576));
    Span4Mux_h I__3223 (
            .O(N__19579),
            .I(N__19573));
    Span4Mux_h I__3222 (
            .O(N__19576),
            .I(N__19570));
    Odrv4 I__3221 (
            .O(N__19573),
            .I(\GENERIC_FIFO_1.n8820 ));
    Odrv4 I__3220 (
            .O(N__19570),
            .I(\GENERIC_FIFO_1.n8820 ));
    InMux I__3219 (
            .O(N__19565),
            .I(N__19560));
    InMux I__3218 (
            .O(N__19564),
            .I(N__19557));
    CascadeMux I__3217 (
            .O(N__19563),
            .I(N__19554));
    LocalMux I__3216 (
            .O(N__19560),
            .I(N__19550));
    LocalMux I__3215 (
            .O(N__19557),
            .I(N__19547));
    InMux I__3214 (
            .O(N__19554),
            .I(N__19544));
    CascadeMux I__3213 (
            .O(N__19553),
            .I(N__19541));
    Span12Mux_v I__3212 (
            .O(N__19550),
            .I(N__19536));
    Span4Mux_v I__3211 (
            .O(N__19547),
            .I(N__19531));
    LocalMux I__3210 (
            .O(N__19544),
            .I(N__19531));
    InMux I__3209 (
            .O(N__19541),
            .I(N__19526));
    InMux I__3208 (
            .O(N__19540),
            .I(N__19526));
    InMux I__3207 (
            .O(N__19539),
            .I(N__19523));
    Odrv12 I__3206 (
            .O(N__19536),
            .I(\GENERIC_FIFO_1.read_pointer_8 ));
    Odrv4 I__3205 (
            .O(N__19531),
            .I(\GENERIC_FIFO_1.read_pointer_8 ));
    LocalMux I__3204 (
            .O(N__19526),
            .I(\GENERIC_FIFO_1.read_pointer_8 ));
    LocalMux I__3203 (
            .O(N__19523),
            .I(\GENERIC_FIFO_1.read_pointer_8 ));
    InMux I__3202 (
            .O(N__19514),
            .I(N__19511));
    LocalMux I__3201 (
            .O(N__19511),
            .I(N__19508));
    Odrv12 I__3200 (
            .O(N__19508),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_0 ));
    SRMux I__3199 (
            .O(N__19505),
            .I(N__19502));
    LocalMux I__3198 (
            .O(N__19502),
            .I(N__19499));
    Span4Mux_h I__3197 (
            .O(N__19499),
            .I(N__19496));
    Odrv4 I__3196 (
            .O(N__19496),
            .I(\Inst_core.Inst_sync.Inst_filter.n4732 ));
    InMux I__3195 (
            .O(N__19493),
            .I(N__19490));
    LocalMux I__3194 (
            .O(N__19490),
            .I(\Inst_core.Inst_sync.Inst_filter.input180Delay_4 ));
    IoInMux I__3193 (
            .O(N__19487),
            .I(N__19484));
    LocalMux I__3192 (
            .O(N__19484),
            .I(N__19481));
    Span4Mux_s0_v I__3191 (
            .O(N__19481),
            .I(N__19477));
    InMux I__3190 (
            .O(N__19480),
            .I(N__19474));
    Odrv4 I__3189 (
            .O(N__19477),
            .I(testcnt_c_0));
    LocalMux I__3188 (
            .O(N__19474),
            .I(testcnt_c_0));
    InMux I__3187 (
            .O(N__19469),
            .I(bfn_6_1_0_));
    InMux I__3186 (
            .O(N__19466),
            .I(N__19463));
    LocalMux I__3185 (
            .O(N__19463),
            .I(N__19460));
    Span4Mux_h I__3184 (
            .O(N__19460),
            .I(N__19457));
    Odrv4 I__3183 (
            .O(N__19457),
            .I(\GENERIC_FIFO_1.n1424 ));
    InMux I__3182 (
            .O(N__19454),
            .I(N__19451));
    LocalMux I__3181 (
            .O(N__19451),
            .I(N__19448));
    Span4Mux_h I__3180 (
            .O(N__19448),
            .I(N__19445));
    Odrv4 I__3179 (
            .O(N__19445),
            .I(\GENERIC_FIFO_1.n1419 ));
    InMux I__3178 (
            .O(N__19442),
            .I(N__19439));
    LocalMux I__3177 (
            .O(N__19439),
            .I(N__19435));
    InMux I__3176 (
            .O(N__19438),
            .I(N__19432));
    Span4Mux_v I__3175 (
            .O(N__19435),
            .I(N__19429));
    LocalMux I__3174 (
            .O(N__19432),
            .I(N__19426));
    Span4Mux_v I__3173 (
            .O(N__19429),
            .I(N__19423));
    Span4Mux_v I__3172 (
            .O(N__19426),
            .I(N__19420));
    Odrv4 I__3171 (
            .O(N__19423),
            .I(\GENERIC_FIFO_1.n8813 ));
    Odrv4 I__3170 (
            .O(N__19420),
            .I(\GENERIC_FIFO_1.n8813 ));
    InMux I__3169 (
            .O(N__19415),
            .I(N__19410));
    InMux I__3168 (
            .O(N__19414),
            .I(N__19407));
    InMux I__3167 (
            .O(N__19413),
            .I(N__19404));
    LocalMux I__3166 (
            .O(N__19410),
            .I(N__19401));
    LocalMux I__3165 (
            .O(N__19407),
            .I(N__19397));
    LocalMux I__3164 (
            .O(N__19404),
            .I(N__19392));
    Span4Mux_h I__3163 (
            .O(N__19401),
            .I(N__19392));
    InMux I__3162 (
            .O(N__19400),
            .I(N__19387));
    Span4Mux_h I__3161 (
            .O(N__19397),
            .I(N__19384));
    Span4Mux_v I__3160 (
            .O(N__19392),
            .I(N__19381));
    InMux I__3159 (
            .O(N__19391),
            .I(N__19378));
    InMux I__3158 (
            .O(N__19390),
            .I(N__19375));
    LocalMux I__3157 (
            .O(N__19387),
            .I(\GENERIC_FIFO_1.read_pointer_1 ));
    Odrv4 I__3156 (
            .O(N__19384),
            .I(\GENERIC_FIFO_1.read_pointer_1 ));
    Odrv4 I__3155 (
            .O(N__19381),
            .I(\GENERIC_FIFO_1.read_pointer_1 ));
    LocalMux I__3154 (
            .O(N__19378),
            .I(\GENERIC_FIFO_1.read_pointer_1 ));
    LocalMux I__3153 (
            .O(N__19375),
            .I(\GENERIC_FIFO_1.read_pointer_1 ));
    InMux I__3152 (
            .O(N__19364),
            .I(N__19361));
    LocalMux I__3151 (
            .O(N__19361),
            .I(N__19357));
    InMux I__3150 (
            .O(N__19360),
            .I(N__19354));
    Span4Mux_v I__3149 (
            .O(N__19357),
            .I(N__19349));
    LocalMux I__3148 (
            .O(N__19354),
            .I(N__19349));
    Span4Mux_h I__3147 (
            .O(N__19349),
            .I(N__19346));
    Odrv4 I__3146 (
            .O(N__19346),
            .I(\GENERIC_FIFO_1.n8814 ));
    InMux I__3145 (
            .O(N__19343),
            .I(N__19339));
    InMux I__3144 (
            .O(N__19342),
            .I(N__19336));
    LocalMux I__3143 (
            .O(N__19339),
            .I(N__19333));
    LocalMux I__3142 (
            .O(N__19336),
            .I(N__19325));
    Span4Mux_h I__3141 (
            .O(N__19333),
            .I(N__19325));
    InMux I__3140 (
            .O(N__19332),
            .I(N__19320));
    InMux I__3139 (
            .O(N__19331),
            .I(N__19320));
    InMux I__3138 (
            .O(N__19330),
            .I(N__19316));
    Span4Mux_v I__3137 (
            .O(N__19325),
            .I(N__19313));
    LocalMux I__3136 (
            .O(N__19320),
            .I(N__19310));
    InMux I__3135 (
            .O(N__19319),
            .I(N__19307));
    LocalMux I__3134 (
            .O(N__19316),
            .I(\GENERIC_FIFO_1.read_pointer_2 ));
    Odrv4 I__3133 (
            .O(N__19313),
            .I(\GENERIC_FIFO_1.read_pointer_2 ));
    Odrv4 I__3132 (
            .O(N__19310),
            .I(\GENERIC_FIFO_1.read_pointer_2 ));
    LocalMux I__3131 (
            .O(N__19307),
            .I(\GENERIC_FIFO_1.read_pointer_2 ));
    InMux I__3130 (
            .O(N__19298),
            .I(N__19295));
    LocalMux I__3129 (
            .O(N__19295),
            .I(N__19292));
    Span4Mux_h I__3128 (
            .O(N__19292),
            .I(N__19289));
    Odrv4 I__3127 (
            .O(N__19289),
            .I(\GENERIC_FIFO_1.n1417 ));
    InMux I__3126 (
            .O(N__19286),
            .I(N__19283));
    LocalMux I__3125 (
            .O(N__19283),
            .I(N__19279));
    InMux I__3124 (
            .O(N__19282),
            .I(N__19276));
    Span4Mux_h I__3123 (
            .O(N__19279),
            .I(N__19273));
    LocalMux I__3122 (
            .O(N__19276),
            .I(N__19270));
    Span4Mux_v I__3121 (
            .O(N__19273),
            .I(N__19267));
    Span4Mux_v I__3120 (
            .O(N__19270),
            .I(N__19264));
    Odrv4 I__3119 (
            .O(N__19267),
            .I(\GENERIC_FIFO_1.n8816 ));
    Odrv4 I__3118 (
            .O(N__19264),
            .I(\GENERIC_FIFO_1.n8816 ));
    InMux I__3117 (
            .O(N__19259),
            .I(N__19255));
    InMux I__3116 (
            .O(N__19258),
            .I(N__19252));
    LocalMux I__3115 (
            .O(N__19255),
            .I(N__19249));
    LocalMux I__3114 (
            .O(N__19252),
            .I(N__19241));
    Span4Mux_h I__3113 (
            .O(N__19249),
            .I(N__19241));
    InMux I__3112 (
            .O(N__19248),
            .I(N__19236));
    InMux I__3111 (
            .O(N__19247),
            .I(N__19236));
    InMux I__3110 (
            .O(N__19246),
            .I(N__19232));
    Span4Mux_v I__3109 (
            .O(N__19241),
            .I(N__19227));
    LocalMux I__3108 (
            .O(N__19236),
            .I(N__19227));
    InMux I__3107 (
            .O(N__19235),
            .I(N__19224));
    LocalMux I__3106 (
            .O(N__19232),
            .I(\GENERIC_FIFO_1.read_pointer_4 ));
    Odrv4 I__3105 (
            .O(N__19227),
            .I(\GENERIC_FIFO_1.read_pointer_4 ));
    LocalMux I__3104 (
            .O(N__19224),
            .I(\GENERIC_FIFO_1.read_pointer_4 ));
    InMux I__3103 (
            .O(N__19217),
            .I(N__19214));
    LocalMux I__3102 (
            .O(N__19214),
            .I(N__19210));
    InMux I__3101 (
            .O(N__19213),
            .I(N__19207));
    Span4Mux_v I__3100 (
            .O(N__19210),
            .I(N__19204));
    LocalMux I__3099 (
            .O(N__19207),
            .I(N__19201));
    Span4Mux_h I__3098 (
            .O(N__19204),
            .I(N__19196));
    Span4Mux_h I__3097 (
            .O(N__19201),
            .I(N__19196));
    Span4Mux_v I__3096 (
            .O(N__19196),
            .I(N__19193));
    Odrv4 I__3095 (
            .O(N__19193),
            .I(\GENERIC_FIFO_1.n8817 ));
    InMux I__3094 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__3093 (
            .O(N__19187),
            .I(N__19183));
    CascadeMux I__3092 (
            .O(N__19186),
            .I(N__19179));
    Span4Mux_v I__3091 (
            .O(N__19183),
            .I(N__19173));
    InMux I__3090 (
            .O(N__19182),
            .I(N__19170));
    InMux I__3089 (
            .O(N__19179),
            .I(N__19165));
    InMux I__3088 (
            .O(N__19178),
            .I(N__19165));
    CascadeMux I__3087 (
            .O(N__19177),
            .I(N__19162));
    InMux I__3086 (
            .O(N__19176),
            .I(N__19159));
    Span4Mux_h I__3085 (
            .O(N__19173),
            .I(N__19156));
    LocalMux I__3084 (
            .O(N__19170),
            .I(N__19151));
    LocalMux I__3083 (
            .O(N__19165),
            .I(N__19151));
    InMux I__3082 (
            .O(N__19162),
            .I(N__19148));
    LocalMux I__3081 (
            .O(N__19159),
            .I(\GENERIC_FIFO_1.read_pointer_5 ));
    Odrv4 I__3080 (
            .O(N__19156),
            .I(\GENERIC_FIFO_1.read_pointer_5 ));
    Odrv4 I__3079 (
            .O(N__19151),
            .I(\GENERIC_FIFO_1.read_pointer_5 ));
    LocalMux I__3078 (
            .O(N__19148),
            .I(\GENERIC_FIFO_1.read_pointer_5 ));
    InMux I__3077 (
            .O(N__19139),
            .I(N__19136));
    LocalMux I__3076 (
            .O(N__19136),
            .I(N__19132));
    InMux I__3075 (
            .O(N__19135),
            .I(N__19129));
    Span4Mux_v I__3074 (
            .O(N__19132),
            .I(N__19124));
    LocalMux I__3073 (
            .O(N__19129),
            .I(N__19124));
    Span4Mux_v I__3072 (
            .O(N__19124),
            .I(N__19121));
    Odrv4 I__3071 (
            .O(N__19121),
            .I(\GENERIC_FIFO_1.n8818 ));
    InMux I__3070 (
            .O(N__19118),
            .I(N__19114));
    CascadeMux I__3069 (
            .O(N__19117),
            .I(N__19111));
    LocalMux I__3068 (
            .O(N__19114),
            .I(N__19106));
    InMux I__3067 (
            .O(N__19111),
            .I(N__19103));
    InMux I__3066 (
            .O(N__19110),
            .I(N__19100));
    InMux I__3065 (
            .O(N__19109),
            .I(N__19095));
    Span12Mux_s4_h I__3064 (
            .O(N__19106),
            .I(N__19092));
    LocalMux I__3063 (
            .O(N__19103),
            .I(N__19087));
    LocalMux I__3062 (
            .O(N__19100),
            .I(N__19087));
    InMux I__3061 (
            .O(N__19099),
            .I(N__19084));
    InMux I__3060 (
            .O(N__19098),
            .I(N__19081));
    LocalMux I__3059 (
            .O(N__19095),
            .I(\GENERIC_FIFO_1.read_pointer_6 ));
    Odrv12 I__3058 (
            .O(N__19092),
            .I(\GENERIC_FIFO_1.read_pointer_6 ));
    Odrv4 I__3057 (
            .O(N__19087),
            .I(\GENERIC_FIFO_1.read_pointer_6 ));
    LocalMux I__3056 (
            .O(N__19084),
            .I(\GENERIC_FIFO_1.read_pointer_6 ));
    LocalMux I__3055 (
            .O(N__19081),
            .I(\GENERIC_FIFO_1.read_pointer_6 ));
    CascadeMux I__3054 (
            .O(N__19070),
            .I(N__19067));
    InMux I__3053 (
            .O(N__19067),
            .I(N__19064));
    LocalMux I__3052 (
            .O(N__19064),
            .I(N__19061));
    Span12Mux_s4_h I__3051 (
            .O(N__19061),
            .I(N__19057));
    InMux I__3050 (
            .O(N__19060),
            .I(N__19054));
    Odrv12 I__3049 (
            .O(N__19057),
            .I(valueRegister_4));
    LocalMux I__3048 (
            .O(N__19054),
            .I(valueRegister_4));
    InMux I__3047 (
            .O(N__19049),
            .I(N__19046));
    LocalMux I__3046 (
            .O(N__19046),
            .I(N__19043));
    Odrv4 I__3045 (
            .O(N__19043),
            .I(\GENERIC_FIFO_1.n1422 ));
    InMux I__3044 (
            .O(N__19040),
            .I(N__19037));
    LocalMux I__3043 (
            .O(N__19037),
            .I(N__19033));
    InMux I__3042 (
            .O(N__19036),
            .I(N__19030));
    Odrv4 I__3041 (
            .O(N__19033),
            .I(valueRegister_7));
    LocalMux I__3040 (
            .O(N__19030),
            .I(valueRegister_7));
    SRMux I__3039 (
            .O(N__19025),
            .I(N__19022));
    LocalMux I__3038 (
            .O(N__19022),
            .I(N__19019));
    Span4Mux_v I__3037 (
            .O(N__19019),
            .I(N__19016));
    Span4Mux_s1_v I__3036 (
            .O(N__19016),
            .I(N__19013));
    Odrv4 I__3035 (
            .O(N__19013),
            .I(\Inst_core.Inst_sync.Inst_filter.n4729 ));
    InMux I__3034 (
            .O(N__19010),
            .I(N__19007));
    LocalMux I__3033 (
            .O(N__19007),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_4 ));
    InMux I__3032 (
            .O(N__19004),
            .I(N__19001));
    LocalMux I__3031 (
            .O(N__19001),
            .I(N__18997));
    InMux I__3030 (
            .O(N__19000),
            .I(N__18994));
    Span4Mux_v I__3029 (
            .O(N__18997),
            .I(N__18989));
    LocalMux I__3028 (
            .O(N__18994),
            .I(N__18989));
    Span4Mux_h I__3027 (
            .O(N__18989),
            .I(N__18986));
    Span4Mux_v I__3026 (
            .O(N__18986),
            .I(N__18983));
    Odrv4 I__3025 (
            .O(N__18983),
            .I(\GENERIC_FIFO_1.n8815 ));
    InMux I__3024 (
            .O(N__18980),
            .I(N__18976));
    InMux I__3023 (
            .O(N__18979),
            .I(N__18973));
    LocalMux I__3022 (
            .O(N__18976),
            .I(N__18970));
    LocalMux I__3021 (
            .O(N__18973),
            .I(N__18964));
    Span4Mux_h I__3020 (
            .O(N__18970),
            .I(N__18964));
    InMux I__3019 (
            .O(N__18969),
            .I(N__18958));
    Span4Mux_v I__3018 (
            .O(N__18964),
            .I(N__18955));
    InMux I__3017 (
            .O(N__18963),
            .I(N__18952));
    InMux I__3016 (
            .O(N__18962),
            .I(N__18949));
    InMux I__3015 (
            .O(N__18961),
            .I(N__18946));
    LocalMux I__3014 (
            .O(N__18958),
            .I(\GENERIC_FIFO_1.read_pointer_3 ));
    Odrv4 I__3013 (
            .O(N__18955),
            .I(\GENERIC_FIFO_1.read_pointer_3 ));
    LocalMux I__3012 (
            .O(N__18952),
            .I(\GENERIC_FIFO_1.read_pointer_3 ));
    LocalMux I__3011 (
            .O(N__18949),
            .I(\GENERIC_FIFO_1.read_pointer_3 ));
    LocalMux I__3010 (
            .O(N__18946),
            .I(\GENERIC_FIFO_1.read_pointer_3 ));
    SRMux I__3009 (
            .O(N__18935),
            .I(N__18932));
    LocalMux I__3008 (
            .O(N__18932),
            .I(N__18929));
    Span12Mux_s6_v I__3007 (
            .O(N__18929),
            .I(N__18926));
    Odrv12 I__3006 (
            .O(N__18926),
            .I(\Inst_core.Inst_sync.Inst_filter.n4731 ));
    InMux I__3005 (
            .O(N__18923),
            .I(N__18919));
    InMux I__3004 (
            .O(N__18922),
            .I(N__18916));
    LocalMux I__3003 (
            .O(N__18919),
            .I(maskRegister_2));
    LocalMux I__3002 (
            .O(N__18916),
            .I(maskRegister_2));
    SRMux I__3001 (
            .O(N__18911),
            .I(N__18908));
    LocalMux I__3000 (
            .O(N__18908),
            .I(N__18905));
    Span4Mux_v I__2999 (
            .O(N__18905),
            .I(N__18902));
    Span4Mux_h I__2998 (
            .O(N__18902),
            .I(N__18899));
    Odrv4 I__2997 (
            .O(N__18899),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4740 ));
    InMux I__2996 (
            .O(N__18896),
            .I(N__18892));
    InMux I__2995 (
            .O(N__18895),
            .I(N__18889));
    LocalMux I__2994 (
            .O(N__18892),
            .I(N__18886));
    LocalMux I__2993 (
            .O(N__18889),
            .I(maskRegister_3));
    Odrv12 I__2992 (
            .O(N__18886),
            .I(maskRegister_3));
    SRMux I__2991 (
            .O(N__18881),
            .I(N__18878));
    LocalMux I__2990 (
            .O(N__18878),
            .I(N__18875));
    Odrv12 I__2989 (
            .O(N__18875),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4741 ));
    InMux I__2988 (
            .O(N__18872),
            .I(N__18868));
    InMux I__2987 (
            .O(N__18871),
            .I(N__18865));
    LocalMux I__2986 (
            .O(N__18868),
            .I(maskRegister_4));
    LocalMux I__2985 (
            .O(N__18865),
            .I(maskRegister_4));
    SRMux I__2984 (
            .O(N__18860),
            .I(N__18857));
    LocalMux I__2983 (
            .O(N__18857),
            .I(N__18854));
    Span4Mux_h I__2982 (
            .O(N__18854),
            .I(N__18851));
    Odrv4 I__2981 (
            .O(N__18851),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4742 ));
    InMux I__2980 (
            .O(N__18848),
            .I(N__18844));
    InMux I__2979 (
            .O(N__18847),
            .I(N__18841));
    LocalMux I__2978 (
            .O(N__18844),
            .I(maskRegister_6));
    LocalMux I__2977 (
            .O(N__18841),
            .I(maskRegister_6));
    SRMux I__2976 (
            .O(N__18836),
            .I(N__18833));
    LocalMux I__2975 (
            .O(N__18833),
            .I(N__18830));
    Span4Mux_v I__2974 (
            .O(N__18830),
            .I(N__18827));
    Odrv4 I__2973 (
            .O(N__18827),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4744 ));
    InMux I__2972 (
            .O(N__18824),
            .I(N__18820));
    InMux I__2971 (
            .O(N__18823),
            .I(N__18817));
    LocalMux I__2970 (
            .O(N__18820),
            .I(maskRegister_7));
    LocalMux I__2969 (
            .O(N__18817),
            .I(maskRegister_7));
    SRMux I__2968 (
            .O(N__18812),
            .I(N__18809));
    LocalMux I__2967 (
            .O(N__18809),
            .I(N__18806));
    Span4Mux_h I__2966 (
            .O(N__18806),
            .I(N__18803));
    Odrv4 I__2965 (
            .O(N__18803),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4745 ));
    InMux I__2964 (
            .O(N__18800),
            .I(N__18794));
    InMux I__2963 (
            .O(N__18799),
            .I(N__18794));
    LocalMux I__2962 (
            .O(N__18794),
            .I(maskRegister_0_adj_1288));
    SRMux I__2961 (
            .O(N__18791),
            .I(N__18788));
    LocalMux I__2960 (
            .O(N__18788),
            .I(N__18785));
    Span4Mux_v I__2959 (
            .O(N__18785),
            .I(N__18782));
    Span4Mux_s1_h I__2958 (
            .O(N__18782),
            .I(N__18779));
    Span4Mux_h I__2957 (
            .O(N__18779),
            .I(N__18776));
    Odrv4 I__2956 (
            .O(N__18776),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4642 ));
    InMux I__2955 (
            .O(N__18773),
            .I(N__18770));
    LocalMux I__2954 (
            .O(N__18770),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_1 ));
    InMux I__2953 (
            .O(N__18767),
            .I(N__18764));
    LocalMux I__2952 (
            .O(N__18764),
            .I(N__18761));
    Odrv4 I__2951 (
            .O(N__18761),
            .I(\Inst_core.Inst_sync.Inst_filter.input360_2 ));
    InMux I__2950 (
            .O(N__18758),
            .I(N__18755));
    LocalMux I__2949 (
            .O(N__18755),
            .I(N__18752));
    Span12Mux_s4_h I__2948 (
            .O(N__18752),
            .I(N__18748));
    InMux I__2947 (
            .O(N__18751),
            .I(N__18745));
    Odrv12 I__2946 (
            .O(N__18748),
            .I(valueRegister_6));
    LocalMux I__2945 (
            .O(N__18745),
            .I(valueRegister_6));
    CascadeMux I__2944 (
            .O(N__18740),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_cascade_ ));
    InMux I__2943 (
            .O(N__18737),
            .I(N__18730));
    InMux I__2942 (
            .O(N__18736),
            .I(N__18730));
    InMux I__2941 (
            .O(N__18735),
            .I(N__18727));
    LocalMux I__2940 (
            .O(N__18730),
            .I(N__18724));
    LocalMux I__2939 (
            .O(N__18727),
            .I(configRegister_23_adj_1339));
    Odrv12 I__2938 (
            .O(N__18724),
            .I(configRegister_23_adj_1339));
    CascadeMux I__2937 (
            .O(N__18719),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9090_cascade_ ));
    SRMux I__2936 (
            .O(N__18716),
            .I(N__18713));
    LocalMux I__2935 (
            .O(N__18713),
            .I(N__18710));
    Odrv4 I__2934 (
            .O(N__18710),
            .I(\Inst_core.Inst_sync.Inst_filter.n4730 ));
    InMux I__2933 (
            .O(N__18707),
            .I(N__18703));
    InMux I__2932 (
            .O(N__18706),
            .I(N__18700));
    LocalMux I__2931 (
            .O(N__18703),
            .I(valueRegister_2));
    LocalMux I__2930 (
            .O(N__18700),
            .I(valueRegister_2));
    CascadeMux I__2929 (
            .O(N__18695),
            .I(N__18692));
    InMux I__2928 (
            .O(N__18692),
            .I(N__18688));
    InMux I__2927 (
            .O(N__18691),
            .I(N__18685));
    LocalMux I__2926 (
            .O(N__18688),
            .I(N__18682));
    LocalMux I__2925 (
            .O(N__18685),
            .I(valueRegister_5));
    Odrv4 I__2924 (
            .O(N__18682),
            .I(valueRegister_5));
    InMux I__2923 (
            .O(N__18677),
            .I(N__18673));
    InMux I__2922 (
            .O(N__18676),
            .I(N__18670));
    LocalMux I__2921 (
            .O(N__18673),
            .I(configRegister_24));
    LocalMux I__2920 (
            .O(N__18670),
            .I(configRegister_24));
    CascadeMux I__2919 (
            .O(N__18665),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9096_cascade_ ));
    CascadeMux I__2918 (
            .O(N__18662),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_cascade_ ));
    InMux I__2917 (
            .O(N__18659),
            .I(N__18654));
    InMux I__2916 (
            .O(N__18658),
            .I(N__18649));
    InMux I__2915 (
            .O(N__18657),
            .I(N__18649));
    LocalMux I__2914 (
            .O(N__18654),
            .I(configRegister_23_adj_1379));
    LocalMux I__2913 (
            .O(N__18649),
            .I(configRegister_23_adj_1379));
    CascadeMux I__2912 (
            .O(N__18644),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9102_cascade_ ));
    InMux I__2911 (
            .O(N__18641),
            .I(N__18637));
    InMux I__2910 (
            .O(N__18640),
            .I(N__18634));
    LocalMux I__2909 (
            .O(N__18637),
            .I(valueRegister_3));
    LocalMux I__2908 (
            .O(N__18634),
            .I(valueRegister_3));
    InMux I__2907 (
            .O(N__18629),
            .I(N__18624));
    InMux I__2906 (
            .O(N__18628),
            .I(N__18619));
    InMux I__2905 (
            .O(N__18627),
            .I(N__18619));
    LocalMux I__2904 (
            .O(N__18624),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3 ));
    LocalMux I__2903 (
            .O(N__18619),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3 ));
    CascadeMux I__2902 (
            .O(N__18614),
            .I(N__18611));
    InMux I__2901 (
            .O(N__18611),
            .I(N__18608));
    LocalMux I__2900 (
            .O(N__18608),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_3 ));
    CascadeMux I__2899 (
            .O(N__18605),
            .I(N__18601));
    CascadeMux I__2898 (
            .O(N__18604),
            .I(N__18598));
    InMux I__2897 (
            .O(N__18601),
            .I(N__18594));
    InMux I__2896 (
            .O(N__18598),
            .I(N__18589));
    InMux I__2895 (
            .O(N__18597),
            .I(N__18589));
    LocalMux I__2894 (
            .O(N__18594),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2 ));
    LocalMux I__2893 (
            .O(N__18589),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2 ));
    InMux I__2892 (
            .O(N__18584),
            .I(N__18581));
    LocalMux I__2891 (
            .O(N__18581),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_2 ));
    CascadeMux I__2890 (
            .O(N__18578),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_cascade_ ));
    CascadeMux I__2889 (
            .O(N__18575),
            .I(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9084_cascade_ ));
    InMux I__2888 (
            .O(N__18572),
            .I(N__18569));
    LocalMux I__2887 (
            .O(N__18569),
            .I(N__18565));
    InMux I__2886 (
            .O(N__18568),
            .I(N__18562));
    Span4Mux_v I__2885 (
            .O(N__18565),
            .I(N__18557));
    LocalMux I__2884 (
            .O(N__18562),
            .I(N__18557));
    Span4Mux_h I__2883 (
            .O(N__18557),
            .I(N__18554));
    Span4Mux_v I__2882 (
            .O(N__18554),
            .I(N__18550));
    InMux I__2881 (
            .O(N__18553),
            .I(N__18547));
    Span4Mux_v I__2880 (
            .O(N__18550),
            .I(N__18544));
    LocalMux I__2879 (
            .O(N__18547),
            .I(\Inst_eia232.Inst_prescaler.counter_1 ));
    Odrv4 I__2878 (
            .O(N__18544),
            .I(\Inst_eia232.Inst_prescaler.counter_1 ));
    InMux I__2877 (
            .O(N__18539),
            .I(N__18536));
    LocalMux I__2876 (
            .O(N__18536),
            .I(N__18532));
    InMux I__2875 (
            .O(N__18535),
            .I(N__18529));
    Span4Mux_h I__2874 (
            .O(N__18532),
            .I(N__18524));
    LocalMux I__2873 (
            .O(N__18529),
            .I(N__18521));
    InMux I__2872 (
            .O(N__18528),
            .I(N__18516));
    InMux I__2871 (
            .O(N__18527),
            .I(N__18516));
    Sp12to4 I__2870 (
            .O(N__18524),
            .I(N__18511));
    Span12Mux_s10_h I__2869 (
            .O(N__18521),
            .I(N__18511));
    LocalMux I__2868 (
            .O(N__18516),
            .I(\Inst_eia232.Inst_prescaler.counter_0 ));
    Odrv12 I__2867 (
            .O(N__18511),
            .I(\Inst_eia232.Inst_prescaler.counter_0 ));
    InMux I__2866 (
            .O(N__18506),
            .I(N__18502));
    InMux I__2865 (
            .O(N__18505),
            .I(N__18499));
    LocalMux I__2864 (
            .O(N__18502),
            .I(N__18496));
    LocalMux I__2863 (
            .O(N__18499),
            .I(N__18493));
    Odrv12 I__2862 (
            .O(N__18496),
            .I(trxClock));
    Odrv12 I__2861 (
            .O(N__18493),
            .I(trxClock));
    CascadeMux I__2860 (
            .O(N__18488),
            .I(N__18485));
    InMux I__2859 (
            .O(N__18485),
            .I(N__18481));
    CascadeMux I__2858 (
            .O(N__18484),
            .I(N__18478));
    LocalMux I__2857 (
            .O(N__18481),
            .I(N__18475));
    InMux I__2856 (
            .O(N__18478),
            .I(N__18472));
    Span4Mux_s2_v I__2855 (
            .O(N__18475),
            .I(N__18465));
    LocalMux I__2854 (
            .O(N__18472),
            .I(N__18465));
    InMux I__2853 (
            .O(N__18471),
            .I(N__18462));
    CascadeMux I__2852 (
            .O(N__18470),
            .I(N__18459));
    Span4Mux_h I__2851 (
            .O(N__18465),
            .I(N__18454));
    LocalMux I__2850 (
            .O(N__18462),
            .I(N__18454));
    InMux I__2849 (
            .O(N__18459),
            .I(N__18451));
    Span4Mux_v I__2848 (
            .O(N__18454),
            .I(N__18446));
    LocalMux I__2847 (
            .O(N__18451),
            .I(N__18446));
    Span4Mux_h I__2846 (
            .O(N__18446),
            .I(N__18443));
    Span4Mux_v I__2845 (
            .O(N__18443),
            .I(N__18440));
    Odrv4 I__2844 (
            .O(N__18440),
            .I(nstate_2__N_139_c_1));
    CascadeMux I__2843 (
            .O(N__18437),
            .I(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_cascade_ ));
    SRMux I__2842 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__2841 (
            .O(N__18431),
            .I(N__18428));
    Span4Mux_s3_v I__2840 (
            .O(N__18428),
            .I(N__18425));
    Span4Mux_v I__2839 (
            .O(N__18425),
            .I(N__18422));
    Span4Mux_v I__2838 (
            .O(N__18422),
            .I(N__18419));
    Odrv4 I__2837 (
            .O(N__18419),
            .I(\Inst_eia232.Inst_prescaler.counter_4__N_38 ));
    InMux I__2836 (
            .O(N__18416),
            .I(N__18409));
    CascadeMux I__2835 (
            .O(N__18415),
            .I(N__18405));
    InMux I__2834 (
            .O(N__18414),
            .I(N__18400));
    InMux I__2833 (
            .O(N__18413),
            .I(N__18400));
    InMux I__2832 (
            .O(N__18412),
            .I(N__18397));
    LocalMux I__2831 (
            .O(N__18409),
            .I(N__18394));
    InMux I__2830 (
            .O(N__18408),
            .I(N__18389));
    InMux I__2829 (
            .O(N__18405),
            .I(N__18389));
    LocalMux I__2828 (
            .O(N__18400),
            .I(\Inst_eia232.Inst_receiver.cmd_4 ));
    LocalMux I__2827 (
            .O(N__18397),
            .I(\Inst_eia232.Inst_receiver.cmd_4 ));
    Odrv4 I__2826 (
            .O(N__18394),
            .I(\Inst_eia232.Inst_receiver.cmd_4 ));
    LocalMux I__2825 (
            .O(N__18389),
            .I(\Inst_eia232.Inst_receiver.cmd_4 ));
    InMux I__2824 (
            .O(N__18380),
            .I(N__18377));
    LocalMux I__2823 (
            .O(N__18377),
            .I(N__18371));
    CascadeMux I__2822 (
            .O(N__18376),
            .I(N__18368));
    CascadeMux I__2821 (
            .O(N__18375),
            .I(N__18365));
    InMux I__2820 (
            .O(N__18374),
            .I(N__18360));
    Span4Mux_h I__2819 (
            .O(N__18371),
            .I(N__18357));
    InMux I__2818 (
            .O(N__18368),
            .I(N__18348));
    InMux I__2817 (
            .O(N__18365),
            .I(N__18348));
    InMux I__2816 (
            .O(N__18364),
            .I(N__18348));
    InMux I__2815 (
            .O(N__18363),
            .I(N__18348));
    LocalMux I__2814 (
            .O(N__18360),
            .I(\Inst_eia232.Inst_receiver.cmd_5 ));
    Odrv4 I__2813 (
            .O(N__18357),
            .I(\Inst_eia232.Inst_receiver.cmd_5 ));
    LocalMux I__2812 (
            .O(N__18348),
            .I(\Inst_eia232.Inst_receiver.cmd_5 ));
    InMux I__2811 (
            .O(N__18341),
            .I(N__18333));
    InMux I__2810 (
            .O(N__18340),
            .I(N__18333));
    InMux I__2809 (
            .O(N__18339),
            .I(N__18328));
    InMux I__2808 (
            .O(N__18338),
            .I(N__18328));
    LocalMux I__2807 (
            .O(N__18333),
            .I(n12));
    LocalMux I__2806 (
            .O(N__18328),
            .I(n12));
    CascadeMux I__2805 (
            .O(N__18323),
            .I(N__18320));
    InMux I__2804 (
            .O(N__18320),
            .I(N__18311));
    InMux I__2803 (
            .O(N__18319),
            .I(N__18311));
    CascadeMux I__2802 (
            .O(N__18318),
            .I(N__18304));
    CascadeMux I__2801 (
            .O(N__18317),
            .I(N__18299));
    CascadeMux I__2800 (
            .O(N__18316),
            .I(N__18296));
    LocalMux I__2799 (
            .O(N__18311),
            .I(N__18290));
    InMux I__2798 (
            .O(N__18310),
            .I(N__18282));
    InMux I__2797 (
            .O(N__18309),
            .I(N__18282));
    InMux I__2796 (
            .O(N__18308),
            .I(N__18282));
    InMux I__2795 (
            .O(N__18307),
            .I(N__18279));
    InMux I__2794 (
            .O(N__18304),
            .I(N__18274));
    InMux I__2793 (
            .O(N__18303),
            .I(N__18274));
    InMux I__2792 (
            .O(N__18302),
            .I(N__18261));
    InMux I__2791 (
            .O(N__18299),
            .I(N__18261));
    InMux I__2790 (
            .O(N__18296),
            .I(N__18261));
    InMux I__2789 (
            .O(N__18295),
            .I(N__18261));
    InMux I__2788 (
            .O(N__18294),
            .I(N__18261));
    InMux I__2787 (
            .O(N__18293),
            .I(N__18261));
    Span4Mux_h I__2786 (
            .O(N__18290),
            .I(N__18258));
    InMux I__2785 (
            .O(N__18289),
            .I(N__18255));
    LocalMux I__2784 (
            .O(N__18282),
            .I(N__18252));
    LocalMux I__2783 (
            .O(N__18279),
            .I(\Inst_eia232.Inst_receiver.cmd_1 ));
    LocalMux I__2782 (
            .O(N__18274),
            .I(\Inst_eia232.Inst_receiver.cmd_1 ));
    LocalMux I__2781 (
            .O(N__18261),
            .I(\Inst_eia232.Inst_receiver.cmd_1 ));
    Odrv4 I__2780 (
            .O(N__18258),
            .I(\Inst_eia232.Inst_receiver.cmd_1 ));
    LocalMux I__2779 (
            .O(N__18255),
            .I(\Inst_eia232.Inst_receiver.cmd_1 ));
    Odrv4 I__2778 (
            .O(N__18252),
            .I(\Inst_eia232.Inst_receiver.cmd_1 ));
    InMux I__2777 (
            .O(N__18239),
            .I(N__18230));
    InMux I__2776 (
            .O(N__18238),
            .I(N__18230));
    InMux I__2775 (
            .O(N__18237),
            .I(N__18230));
    LocalMux I__2774 (
            .O(N__18230),
            .I(N__18222));
    InMux I__2773 (
            .O(N__18229),
            .I(N__18211));
    InMux I__2772 (
            .O(N__18228),
            .I(N__18211));
    InMux I__2771 (
            .O(N__18227),
            .I(N__18211));
    InMux I__2770 (
            .O(N__18226),
            .I(N__18211));
    InMux I__2769 (
            .O(N__18225),
            .I(N__18211));
    Span4Mux_v I__2768 (
            .O(N__18222),
            .I(N__18208));
    LocalMux I__2767 (
            .O(N__18211),
            .I(\Inst_eia232.Inst_receiver.n3718 ));
    Odrv4 I__2766 (
            .O(N__18208),
            .I(\Inst_eia232.Inst_receiver.n3718 ));
    CascadeMux I__2765 (
            .O(N__18203),
            .I(N__18195));
    CascadeMux I__2764 (
            .O(N__18202),
            .I(N__18190));
    CascadeMux I__2763 (
            .O(N__18201),
            .I(N__18186));
    CascadeMux I__2762 (
            .O(N__18200),
            .I(N__18183));
    CascadeMux I__2761 (
            .O(N__18199),
            .I(N__18180));
    CascadeMux I__2760 (
            .O(N__18198),
            .I(N__18174));
    InMux I__2759 (
            .O(N__18195),
            .I(N__18166));
    InMux I__2758 (
            .O(N__18194),
            .I(N__18166));
    InMux I__2757 (
            .O(N__18193),
            .I(N__18166));
    InMux I__2756 (
            .O(N__18190),
            .I(N__18163));
    InMux I__2755 (
            .O(N__18189),
            .I(N__18148));
    InMux I__2754 (
            .O(N__18186),
            .I(N__18148));
    InMux I__2753 (
            .O(N__18183),
            .I(N__18148));
    InMux I__2752 (
            .O(N__18180),
            .I(N__18148));
    InMux I__2751 (
            .O(N__18179),
            .I(N__18148));
    InMux I__2750 (
            .O(N__18178),
            .I(N__18148));
    InMux I__2749 (
            .O(N__18177),
            .I(N__18148));
    InMux I__2748 (
            .O(N__18174),
            .I(N__18143));
    InMux I__2747 (
            .O(N__18173),
            .I(N__18143));
    LocalMux I__2746 (
            .O(N__18166),
            .I(N__18140));
    LocalMux I__2745 (
            .O(N__18163),
            .I(\Inst_eia232.Inst_receiver.cmd_2 ));
    LocalMux I__2744 (
            .O(N__18148),
            .I(\Inst_eia232.Inst_receiver.cmd_2 ));
    LocalMux I__2743 (
            .O(N__18143),
            .I(\Inst_eia232.Inst_receiver.cmd_2 ));
    Odrv4 I__2742 (
            .O(N__18140),
            .I(\Inst_eia232.Inst_receiver.cmd_2 ));
    InMux I__2741 (
            .O(N__18131),
            .I(N__18115));
    InMux I__2740 (
            .O(N__18130),
            .I(N__18115));
    InMux I__2739 (
            .O(N__18129),
            .I(N__18115));
    InMux I__2738 (
            .O(N__18128),
            .I(N__18098));
    InMux I__2737 (
            .O(N__18127),
            .I(N__18098));
    InMux I__2736 (
            .O(N__18126),
            .I(N__18098));
    InMux I__2735 (
            .O(N__18125),
            .I(N__18098));
    InMux I__2734 (
            .O(N__18124),
            .I(N__18098));
    InMux I__2733 (
            .O(N__18123),
            .I(N__18098));
    InMux I__2732 (
            .O(N__18122),
            .I(N__18098));
    LocalMux I__2731 (
            .O(N__18115),
            .I(N__18095));
    InMux I__2730 (
            .O(N__18114),
            .I(N__18090));
    InMux I__2729 (
            .O(N__18113),
            .I(N__18090));
    LocalMux I__2728 (
            .O(N__18098),
            .I(\Inst_eia232.Inst_receiver.cmd_0 ));
    Odrv4 I__2727 (
            .O(N__18095),
            .I(\Inst_eia232.Inst_receiver.cmd_0 ));
    LocalMux I__2726 (
            .O(N__18090),
            .I(\Inst_eia232.Inst_receiver.cmd_0 ));
    CascadeMux I__2725 (
            .O(N__18083),
            .I(N__18076));
    CascadeMux I__2724 (
            .O(N__18082),
            .I(N__18070));
    CascadeMux I__2723 (
            .O(N__18081),
            .I(N__18066));
    InMux I__2722 (
            .O(N__18080),
            .I(N__18061));
    InMux I__2721 (
            .O(N__18079),
            .I(N__18061));
    InMux I__2720 (
            .O(N__18076),
            .I(N__18042));
    InMux I__2719 (
            .O(N__18075),
            .I(N__18042));
    InMux I__2718 (
            .O(N__18074),
            .I(N__18042));
    InMux I__2717 (
            .O(N__18073),
            .I(N__18042));
    InMux I__2716 (
            .O(N__18070),
            .I(N__18042));
    InMux I__2715 (
            .O(N__18069),
            .I(N__18042));
    InMux I__2714 (
            .O(N__18066),
            .I(N__18042));
    LocalMux I__2713 (
            .O(N__18061),
            .I(N__18039));
    InMux I__2712 (
            .O(N__18060),
            .I(N__18036));
    InMux I__2711 (
            .O(N__18059),
            .I(N__18029));
    InMux I__2710 (
            .O(N__18058),
            .I(N__18029));
    InMux I__2709 (
            .O(N__18057),
            .I(N__18029));
    LocalMux I__2708 (
            .O(N__18042),
            .I(N__18024));
    Span4Mux_h I__2707 (
            .O(N__18039),
            .I(N__18024));
    LocalMux I__2706 (
            .O(N__18036),
            .I(\Inst_eia232.Inst_receiver.cmd_3 ));
    LocalMux I__2705 (
            .O(N__18029),
            .I(\Inst_eia232.Inst_receiver.cmd_3 ));
    Odrv4 I__2704 (
            .O(N__18024),
            .I(\Inst_eia232.Inst_receiver.cmd_3 ));
    CascadeMux I__2703 (
            .O(N__18017),
            .I(N__18013));
    InMux I__2702 (
            .O(N__18016),
            .I(N__18010));
    InMux I__2701 (
            .O(N__18013),
            .I(N__18003));
    LocalMux I__2700 (
            .O(N__18010),
            .I(N__18000));
    InMux I__2699 (
            .O(N__18009),
            .I(N__17991));
    InMux I__2698 (
            .O(N__18008),
            .I(N__17991));
    InMux I__2697 (
            .O(N__18007),
            .I(N__17991));
    InMux I__2696 (
            .O(N__18006),
            .I(N__17991));
    LocalMux I__2695 (
            .O(N__18003),
            .I(\Inst_eia232.Inst_receiver.n69 ));
    Odrv4 I__2694 (
            .O(N__18000),
            .I(\Inst_eia232.Inst_receiver.n69 ));
    LocalMux I__2693 (
            .O(N__17991),
            .I(\Inst_eia232.Inst_receiver.n69 ));
    InMux I__2692 (
            .O(N__17984),
            .I(N__17977));
    InMux I__2691 (
            .O(N__17983),
            .I(N__17977));
    CascadeMux I__2690 (
            .O(N__17982),
            .I(N__17972));
    LocalMux I__2689 (
            .O(N__17977),
            .I(N__17968));
    InMux I__2688 (
            .O(N__17976),
            .I(N__17962));
    InMux I__2687 (
            .O(N__17975),
            .I(N__17959));
    InMux I__2686 (
            .O(N__17972),
            .I(N__17954));
    InMux I__2685 (
            .O(N__17971),
            .I(N__17954));
    Span4Mux_h I__2684 (
            .O(N__17968),
            .I(N__17951));
    CascadeMux I__2683 (
            .O(N__17967),
            .I(N__17947));
    CascadeMux I__2682 (
            .O(N__17966),
            .I(N__17943));
    CascadeMux I__2681 (
            .O(N__17965),
            .I(N__17939));
    LocalMux I__2680 (
            .O(N__17962),
            .I(N__17932));
    LocalMux I__2679 (
            .O(N__17959),
            .I(N__17925));
    LocalMux I__2678 (
            .O(N__17954),
            .I(N__17925));
    Span4Mux_v I__2677 (
            .O(N__17951),
            .I(N__17925));
    InMux I__2676 (
            .O(N__17950),
            .I(N__17922));
    InMux I__2675 (
            .O(N__17947),
            .I(N__17911));
    InMux I__2674 (
            .O(N__17946),
            .I(N__17911));
    InMux I__2673 (
            .O(N__17943),
            .I(N__17911));
    InMux I__2672 (
            .O(N__17942),
            .I(N__17911));
    InMux I__2671 (
            .O(N__17939),
            .I(N__17911));
    InMux I__2670 (
            .O(N__17938),
            .I(N__17904));
    InMux I__2669 (
            .O(N__17937),
            .I(N__17904));
    InMux I__2668 (
            .O(N__17936),
            .I(N__17904));
    InMux I__2667 (
            .O(N__17935),
            .I(N__17901));
    Span4Mux_h I__2666 (
            .O(N__17932),
            .I(N__17896));
    Span4Mux_v I__2665 (
            .O(N__17925),
            .I(N__17896));
    LocalMux I__2664 (
            .O(N__17922),
            .I(\Inst_eia232.state_1 ));
    LocalMux I__2663 (
            .O(N__17911),
            .I(\Inst_eia232.state_1 ));
    LocalMux I__2662 (
            .O(N__17904),
            .I(\Inst_eia232.state_1 ));
    LocalMux I__2661 (
            .O(N__17901),
            .I(\Inst_eia232.state_1 ));
    Odrv4 I__2660 (
            .O(N__17896),
            .I(\Inst_eia232.state_1 ));
    InMux I__2659 (
            .O(N__17885),
            .I(N__17876));
    InMux I__2658 (
            .O(N__17884),
            .I(N__17876));
    InMux I__2657 (
            .O(N__17883),
            .I(N__17873));
    InMux I__2656 (
            .O(N__17882),
            .I(N__17870));
    InMux I__2655 (
            .O(N__17881),
            .I(N__17867));
    LocalMux I__2654 (
            .O(N__17876),
            .I(N__17864));
    LocalMux I__2653 (
            .O(N__17873),
            .I(N__17847));
    LocalMux I__2652 (
            .O(N__17870),
            .I(N__17847));
    LocalMux I__2651 (
            .O(N__17867),
            .I(N__17847));
    Span4Mux_v I__2650 (
            .O(N__17864),
            .I(N__17847));
    CascadeMux I__2649 (
            .O(N__17863),
            .I(N__17843));
    InMux I__2648 (
            .O(N__17862),
            .I(N__17838));
    InMux I__2647 (
            .O(N__17861),
            .I(N__17835));
    InMux I__2646 (
            .O(N__17860),
            .I(N__17824));
    InMux I__2645 (
            .O(N__17859),
            .I(N__17824));
    InMux I__2644 (
            .O(N__17858),
            .I(N__17824));
    InMux I__2643 (
            .O(N__17857),
            .I(N__17824));
    InMux I__2642 (
            .O(N__17856),
            .I(N__17824));
    Span4Mux_v I__2641 (
            .O(N__17847),
            .I(N__17821));
    InMux I__2640 (
            .O(N__17846),
            .I(N__17812));
    InMux I__2639 (
            .O(N__17843),
            .I(N__17812));
    InMux I__2638 (
            .O(N__17842),
            .I(N__17812));
    InMux I__2637 (
            .O(N__17841),
            .I(N__17812));
    LocalMux I__2636 (
            .O(N__17838),
            .I(\Inst_eia232.state_2 ));
    LocalMux I__2635 (
            .O(N__17835),
            .I(\Inst_eia232.state_2 ));
    LocalMux I__2634 (
            .O(N__17824),
            .I(\Inst_eia232.state_2 ));
    Odrv4 I__2633 (
            .O(N__17821),
            .I(\Inst_eia232.state_2 ));
    LocalMux I__2632 (
            .O(N__17812),
            .I(\Inst_eia232.state_2 ));
    CascadeMux I__2631 (
            .O(N__17801),
            .I(\Inst_eia232.Inst_receiver.n7_cascade_ ));
    InMux I__2630 (
            .O(N__17798),
            .I(N__17788));
    InMux I__2629 (
            .O(N__17797),
            .I(N__17788));
    InMux I__2628 (
            .O(N__17796),
            .I(N__17779));
    InMux I__2627 (
            .O(N__17795),
            .I(N__17779));
    InMux I__2626 (
            .O(N__17794),
            .I(N__17779));
    InMux I__2625 (
            .O(N__17793),
            .I(N__17779));
    LocalMux I__2624 (
            .O(N__17788),
            .I(\Inst_eia232.Inst_receiver.counter_1 ));
    LocalMux I__2623 (
            .O(N__17779),
            .I(\Inst_eia232.Inst_receiver.counter_1 ));
    InMux I__2622 (
            .O(N__17774),
            .I(N__17763));
    InMux I__2621 (
            .O(N__17773),
            .I(N__17763));
    InMux I__2620 (
            .O(N__17772),
            .I(N__17752));
    InMux I__2619 (
            .O(N__17771),
            .I(N__17752));
    InMux I__2618 (
            .O(N__17770),
            .I(N__17752));
    InMux I__2617 (
            .O(N__17769),
            .I(N__17752));
    InMux I__2616 (
            .O(N__17768),
            .I(N__17752));
    LocalMux I__2615 (
            .O(N__17763),
            .I(\Inst_eia232.Inst_receiver.counter_0 ));
    LocalMux I__2614 (
            .O(N__17752),
            .I(\Inst_eia232.Inst_receiver.counter_0 ));
    CascadeMux I__2613 (
            .O(N__17747),
            .I(N__17741));
    InMux I__2612 (
            .O(N__17746),
            .I(N__17735));
    InMux I__2611 (
            .O(N__17745),
            .I(N__17735));
    InMux I__2610 (
            .O(N__17744),
            .I(N__17728));
    InMux I__2609 (
            .O(N__17741),
            .I(N__17728));
    InMux I__2608 (
            .O(N__17740),
            .I(N__17728));
    LocalMux I__2607 (
            .O(N__17735),
            .I(\Inst_eia232.Inst_receiver.counter_2 ));
    LocalMux I__2606 (
            .O(N__17728),
            .I(\Inst_eia232.Inst_receiver.counter_2 ));
    InMux I__2605 (
            .O(N__17723),
            .I(N__17720));
    LocalMux I__2604 (
            .O(N__17720),
            .I(\Inst_eia232.Inst_receiver.n7777 ));
    SRMux I__2603 (
            .O(N__17717),
            .I(N__17714));
    LocalMux I__2602 (
            .O(N__17714),
            .I(N__17711));
    Span4Mux_s0_v I__2601 (
            .O(N__17711),
            .I(N__17708));
    Odrv4 I__2600 (
            .O(N__17708),
            .I(\Inst_eia232.Inst_receiver.n3202 ));
    InMux I__2599 (
            .O(N__17705),
            .I(N__17702));
    LocalMux I__2598 (
            .O(N__17702),
            .I(N__17699));
    Odrv12 I__2597 (
            .O(N__17699),
            .I(\Inst_eia232.Inst_receiver.n1_adj_1266 ));
    InMux I__2596 (
            .O(N__17696),
            .I(N__17687));
    InMux I__2595 (
            .O(N__17695),
            .I(N__17687));
    InMux I__2594 (
            .O(N__17694),
            .I(N__17680));
    InMux I__2593 (
            .O(N__17693),
            .I(N__17680));
    InMux I__2592 (
            .O(N__17692),
            .I(N__17680));
    LocalMux I__2591 (
            .O(N__17687),
            .I(N__17677));
    LocalMux I__2590 (
            .O(N__17680),
            .I(N__17668));
    Span4Mux_v I__2589 (
            .O(N__17677),
            .I(N__17668));
    CascadeMux I__2588 (
            .O(N__17676),
            .I(N__17665));
    CascadeMux I__2587 (
            .O(N__17675),
            .I(N__17658));
    InMux I__2586 (
            .O(N__17674),
            .I(N__17650));
    InMux I__2585 (
            .O(N__17673),
            .I(N__17647));
    Span4Mux_v I__2584 (
            .O(N__17668),
            .I(N__17644));
    InMux I__2583 (
            .O(N__17665),
            .I(N__17633));
    InMux I__2582 (
            .O(N__17664),
            .I(N__17633));
    InMux I__2581 (
            .O(N__17663),
            .I(N__17633));
    InMux I__2580 (
            .O(N__17662),
            .I(N__17633));
    InMux I__2579 (
            .O(N__17661),
            .I(N__17633));
    InMux I__2578 (
            .O(N__17658),
            .I(N__17630));
    InMux I__2577 (
            .O(N__17657),
            .I(N__17619));
    InMux I__2576 (
            .O(N__17656),
            .I(N__17619));
    InMux I__2575 (
            .O(N__17655),
            .I(N__17619));
    InMux I__2574 (
            .O(N__17654),
            .I(N__17619));
    InMux I__2573 (
            .O(N__17653),
            .I(N__17619));
    LocalMux I__2572 (
            .O(N__17650),
            .I(\Inst_eia232.state_0 ));
    LocalMux I__2571 (
            .O(N__17647),
            .I(\Inst_eia232.state_0 ));
    Odrv4 I__2570 (
            .O(N__17644),
            .I(\Inst_eia232.state_0 ));
    LocalMux I__2569 (
            .O(N__17633),
            .I(\Inst_eia232.state_0 ));
    LocalMux I__2568 (
            .O(N__17630),
            .I(\Inst_eia232.state_0 ));
    LocalMux I__2567 (
            .O(N__17619),
            .I(\Inst_eia232.state_0 ));
    InMux I__2566 (
            .O(N__17606),
            .I(N__17599));
    InMux I__2565 (
            .O(N__17605),
            .I(N__17592));
    InMux I__2564 (
            .O(N__17604),
            .I(N__17592));
    InMux I__2563 (
            .O(N__17603),
            .I(N__17592));
    InMux I__2562 (
            .O(N__17602),
            .I(N__17589));
    LocalMux I__2561 (
            .O(N__17599),
            .I(N__17584));
    LocalMux I__2560 (
            .O(N__17592),
            .I(N__17584));
    LocalMux I__2559 (
            .O(N__17589),
            .I(\Inst_eia232.Inst_receiver.nstate_2_N_133_1 ));
    Odrv4 I__2558 (
            .O(N__17584),
            .I(\Inst_eia232.Inst_receiver.nstate_2_N_133_1 ));
    InMux I__2557 (
            .O(N__17579),
            .I(N__17576));
    LocalMux I__2556 (
            .O(N__17576),
            .I(N__17573));
    Odrv12 I__2555 (
            .O(N__17573),
            .I(\Inst_eia232.Inst_receiver.n8826 ));
    CascadeMux I__2554 (
            .O(N__17570),
            .I(\Inst_eia232.Inst_receiver.n3504_cascade_ ));
    CEMux I__2553 (
            .O(N__17567),
            .I(N__17564));
    LocalMux I__2552 (
            .O(N__17564),
            .I(N__17561));
    Span4Mux_v I__2551 (
            .O(N__17561),
            .I(N__17558));
    Span4Mux_s0_v I__2550 (
            .O(N__17558),
            .I(N__17555));
    Odrv4 I__2549 (
            .O(N__17555),
            .I(\Inst_eia232.Inst_receiver.n3676 ));
    SRMux I__2548 (
            .O(N__17552),
            .I(N__17549));
    LocalMux I__2547 (
            .O(N__17549),
            .I(N__17546));
    Span4Mux_v I__2546 (
            .O(N__17546),
            .I(N__17543));
    Odrv4 I__2545 (
            .O(N__17543),
            .I(\Inst_eia232.Inst_receiver.n4767 ));
    InMux I__2544 (
            .O(N__17540),
            .I(N__17537));
    LocalMux I__2543 (
            .O(N__17537),
            .I(\Inst_eia232.Inst_receiver.n3504 ));
    InMux I__2542 (
            .O(N__17534),
            .I(N__17528));
    InMux I__2541 (
            .O(N__17533),
            .I(N__17528));
    LocalMux I__2540 (
            .O(N__17528),
            .I(N__17525));
    Odrv4 I__2539 (
            .O(N__17525),
            .I(\Inst_eia232.Inst_receiver.n5 ));
    InMux I__2538 (
            .O(N__17522),
            .I(N__17515));
    InMux I__2537 (
            .O(N__17521),
            .I(N__17515));
    InMux I__2536 (
            .O(N__17520),
            .I(N__17512));
    LocalMux I__2535 (
            .O(N__17515),
            .I(\Inst_eia232.Inst_receiver.n75 ));
    LocalMux I__2534 (
            .O(N__17512),
            .I(\Inst_eia232.Inst_receiver.n75 ));
    CascadeMux I__2533 (
            .O(N__17507),
            .I(N__17504));
    InMux I__2532 (
            .O(N__17504),
            .I(N__17498));
    InMux I__2531 (
            .O(N__17503),
            .I(N__17498));
    LocalMux I__2530 (
            .O(N__17498),
            .I(\Inst_eia232.Inst_receiver.n14 ));
    SRMux I__2529 (
            .O(N__17495),
            .I(N__17491));
    SRMux I__2528 (
            .O(N__17494),
            .I(N__17488));
    LocalMux I__2527 (
            .O(N__17491),
            .I(N__17483));
    LocalMux I__2526 (
            .O(N__17488),
            .I(N__17480));
    SRMux I__2525 (
            .O(N__17487),
            .I(N__17477));
    SRMux I__2524 (
            .O(N__17486),
            .I(N__17474));
    Span4Mux_v I__2523 (
            .O(N__17483),
            .I(N__17471));
    Span4Mux_v I__2522 (
            .O(N__17480),
            .I(N__17464));
    LocalMux I__2521 (
            .O(N__17477),
            .I(N__17464));
    LocalMux I__2520 (
            .O(N__17474),
            .I(N__17464));
    Odrv4 I__2519 (
            .O(N__17471),
            .I(n1917));
    Odrv4 I__2518 (
            .O(N__17464),
            .I(n1917));
    InMux I__2517 (
            .O(N__17459),
            .I(N__17449));
    InMux I__2516 (
            .O(N__17458),
            .I(N__17449));
    InMux I__2515 (
            .O(N__17457),
            .I(N__17449));
    InMux I__2514 (
            .O(N__17456),
            .I(N__17446));
    LocalMux I__2513 (
            .O(N__17449),
            .I(\Inst_eia232.Inst_receiver.counter_4 ));
    LocalMux I__2512 (
            .O(N__17446),
            .I(\Inst_eia232.Inst_receiver.counter_4 ));
    CascadeMux I__2511 (
            .O(N__17441),
            .I(N__17436));
    InMux I__2510 (
            .O(N__17440),
            .I(N__17431));
    InMux I__2509 (
            .O(N__17439),
            .I(N__17428));
    InMux I__2508 (
            .O(N__17436),
            .I(N__17421));
    InMux I__2507 (
            .O(N__17435),
            .I(N__17421));
    InMux I__2506 (
            .O(N__17434),
            .I(N__17421));
    LocalMux I__2505 (
            .O(N__17431),
            .I(\Inst_eia232.Inst_receiver.counter_3 ));
    LocalMux I__2504 (
            .O(N__17428),
            .I(\Inst_eia232.Inst_receiver.counter_3 ));
    LocalMux I__2503 (
            .O(N__17421),
            .I(\Inst_eia232.Inst_receiver.counter_3 ));
    InMux I__2502 (
            .O(N__17414),
            .I(N__17409));
    InMux I__2501 (
            .O(N__17413),
            .I(N__17404));
    InMux I__2500 (
            .O(N__17412),
            .I(N__17404));
    LocalMux I__2499 (
            .O(N__17409),
            .I(\Inst_eia232.Inst_receiver.n5504 ));
    LocalMux I__2498 (
            .O(N__17404),
            .I(\Inst_eia232.Inst_receiver.n5504 ));
    CascadeMux I__2497 (
            .O(N__17399),
            .I(\Inst_eia232.Inst_receiver.n8782_cascade_ ));
    InMux I__2496 (
            .O(N__17396),
            .I(N__17390));
    InMux I__2495 (
            .O(N__17395),
            .I(N__17390));
    LocalMux I__2494 (
            .O(N__17390),
            .I(\Inst_eia232.Inst_receiver.n6_adj_1267 ));
    CascadeMux I__2493 (
            .O(N__17387),
            .I(\Inst_eia232.Inst_receiver.n3_cascade_ ));
    InMux I__2492 (
            .O(N__17384),
            .I(N__17381));
    LocalMux I__2491 (
            .O(N__17381),
            .I(\Inst_eia232.Inst_receiver.n5505 ));
    CascadeMux I__2490 (
            .O(N__17378),
            .I(\Inst_eia232.Inst_receiver.n8755_cascade_ ));
    CascadeMux I__2489 (
            .O(N__17375),
            .I(\Inst_eia232.Inst_receiver.n9123_cascade_ ));
    InMux I__2488 (
            .O(N__17372),
            .I(N__17369));
    LocalMux I__2487 (
            .O(N__17369),
            .I(executePrev));
    InMux I__2486 (
            .O(N__17366),
            .I(N__17363));
    LocalMux I__2485 (
            .O(N__17363),
            .I(\Inst_eia232.Inst_receiver.n8784 ));
    CascadeMux I__2484 (
            .O(N__17360),
            .I(\Inst_eia232.Inst_receiver.n6_cascade_ ));
    CascadeMux I__2483 (
            .O(N__17357),
            .I(\Inst_eia232.Inst_receiver.n8_cascade_ ));
    SRMux I__2482 (
            .O(N__17354),
            .I(N__17351));
    LocalMux I__2481 (
            .O(N__17351),
            .I(N__17346));
    SRMux I__2480 (
            .O(N__17350),
            .I(N__17343));
    InMux I__2479 (
            .O(N__17349),
            .I(N__17340));
    Span4Mux_v I__2478 (
            .O(N__17346),
            .I(N__17335));
    LocalMux I__2477 (
            .O(N__17343),
            .I(N__17335));
    LocalMux I__2476 (
            .O(N__17340),
            .I(N__17332));
    Span4Mux_v I__2475 (
            .O(N__17335),
            .I(N__17329));
    Odrv12 I__2474 (
            .O(N__17332),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2473 (
            .O(N__17329),
            .I(CONSTANT_ONE_NET));
    InMux I__2472 (
            .O(N__17324),
            .I(N__17321));
    LocalMux I__2471 (
            .O(N__17321),
            .I(\GENERIC_FIFO_1.n1388 ));
    CascadeMux I__2470 (
            .O(N__17318),
            .I(N__17315));
    InMux I__2469 (
            .O(N__17315),
            .I(N__17312));
    LocalMux I__2468 (
            .O(N__17312),
            .I(N__17309));
    Odrv4 I__2467 (
            .O(N__17309),
            .I(\GENERIC_FIFO_1.n1373 ));
    InMux I__2466 (
            .O(N__17306),
            .I(N__17303));
    LocalMux I__2465 (
            .O(N__17303),
            .I(N__17300));
    Span4Mux_s3_h I__2464 (
            .O(N__17300),
            .I(N__17297));
    Span4Mux_v I__2463 (
            .O(N__17297),
            .I(N__17294));
    Odrv4 I__2462 (
            .O(N__17294),
            .I(\GENERIC_FIFO_1.n8630 ));
    InMux I__2461 (
            .O(N__17291),
            .I(bfn_4_16_0_));
    CascadeMux I__2460 (
            .O(N__17288),
            .I(N__17285));
    InMux I__2459 (
            .O(N__17285),
            .I(N__17282));
    LocalMux I__2458 (
            .O(N__17282),
            .I(N__17279));
    Odrv4 I__2457 (
            .O(N__17279),
            .I(\GENERIC_FIFO_1.n1372 ));
    InMux I__2456 (
            .O(N__17276),
            .I(\GENERIC_FIFO_1.n7945 ));
    InMux I__2455 (
            .O(N__17273),
            .I(N__17270));
    LocalMux I__2454 (
            .O(N__17270),
            .I(\GENERIC_FIFO_1.n1383 ));
    CascadeMux I__2453 (
            .O(N__17267),
            .I(N__17264));
    InMux I__2452 (
            .O(N__17264),
            .I(N__17261));
    LocalMux I__2451 (
            .O(N__17261),
            .I(N__17258));
    Odrv4 I__2450 (
            .O(N__17258),
            .I(\GENERIC_FIFO_1.n1371 ));
    InMux I__2449 (
            .O(N__17255),
            .I(N__17252));
    LocalMux I__2448 (
            .O(N__17252),
            .I(N__17249));
    Span4Mux_v I__2447 (
            .O(N__17249),
            .I(N__17246));
    Span4Mux_v I__2446 (
            .O(N__17246),
            .I(N__17243));
    Odrv4 I__2445 (
            .O(N__17243),
            .I(\GENERIC_FIFO_1.n8638 ));
    InMux I__2444 (
            .O(N__17240),
            .I(\GENERIC_FIFO_1.n7946 ));
    InMux I__2443 (
            .O(N__17237),
            .I(\GENERIC_FIFO_1.n1392 ));
    InMux I__2442 (
            .O(N__17234),
            .I(N__17230));
    InMux I__2441 (
            .O(N__17233),
            .I(N__17226));
    LocalMux I__2440 (
            .O(N__17230),
            .I(N__17223));
    InMux I__2439 (
            .O(N__17229),
            .I(N__17220));
    LocalMux I__2438 (
            .O(N__17226),
            .I(N__17217));
    Span4Mux_v I__2437 (
            .O(N__17223),
            .I(N__17212));
    LocalMux I__2436 (
            .O(N__17220),
            .I(N__17212));
    Span4Mux_s3_h I__2435 (
            .O(N__17217),
            .I(N__17209));
    Span4Mux_v I__2434 (
            .O(N__17212),
            .I(N__17206));
    Odrv4 I__2433 (
            .O(N__17209),
            .I(\GENERIC_FIFO_1.n1392_THRU_CO ));
    Odrv4 I__2432 (
            .O(N__17206),
            .I(\GENERIC_FIFO_1.n1392_THRU_CO ));
    InMux I__2431 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__2430 (
            .O(N__17198),
            .I(N__17195));
    Span4Mux_s3_v I__2429 (
            .O(N__17195),
            .I(N__17191));
    InMux I__2428 (
            .O(N__17194),
            .I(N__17188));
    Span4Mux_v I__2427 (
            .O(N__17191),
            .I(N__17185));
    LocalMux I__2426 (
            .O(N__17188),
            .I(N__17182));
    Odrv4 I__2425 (
            .O(N__17185),
            .I(\GENERIC_FIFO_1.n8821 ));
    Odrv12 I__2424 (
            .O(N__17182),
            .I(\GENERIC_FIFO_1.n8821 ));
    InMux I__2423 (
            .O(N__17177),
            .I(N__17173));
    InMux I__2422 (
            .O(N__17176),
            .I(N__17169));
    LocalMux I__2421 (
            .O(N__17173),
            .I(N__17166));
    CascadeMux I__2420 (
            .O(N__17172),
            .I(N__17163));
    LocalMux I__2419 (
            .O(N__17169),
            .I(N__17158));
    Span4Mux_v I__2418 (
            .O(N__17166),
            .I(N__17158));
    InMux I__2417 (
            .O(N__17163),
            .I(N__17155));
    Span4Mux_v I__2416 (
            .O(N__17158),
            .I(N__17149));
    LocalMux I__2415 (
            .O(N__17155),
            .I(N__17146));
    InMux I__2414 (
            .O(N__17154),
            .I(N__17139));
    InMux I__2413 (
            .O(N__17153),
            .I(N__17139));
    InMux I__2412 (
            .O(N__17152),
            .I(N__17139));
    Odrv4 I__2411 (
            .O(N__17149),
            .I(\GENERIC_FIFO_1.read_pointer_9 ));
    Odrv4 I__2410 (
            .O(N__17146),
            .I(\GENERIC_FIFO_1.read_pointer_9 ));
    LocalMux I__2409 (
            .O(N__17139),
            .I(\GENERIC_FIFO_1.read_pointer_9 ));
    InMux I__2408 (
            .O(N__17132),
            .I(N__17129));
    LocalMux I__2407 (
            .O(N__17129),
            .I(N__17126));
    Span4Mux_s3_h I__2406 (
            .O(N__17126),
            .I(N__17123));
    Odrv4 I__2405 (
            .O(N__17123),
            .I(\GENERIC_FIFO_1.n1416 ));
    CascadeMux I__2404 (
            .O(N__17120),
            .I(N__17117));
    CascadeBuf I__2403 (
            .O(N__17117),
            .I(N__17112));
    InMux I__2402 (
            .O(N__17116),
            .I(N__17109));
    InMux I__2401 (
            .O(N__17115),
            .I(N__17106));
    CascadeMux I__2400 (
            .O(N__17112),
            .I(N__17103));
    LocalMux I__2399 (
            .O(N__17109),
            .I(N__17098));
    LocalMux I__2398 (
            .O(N__17106),
            .I(N__17095));
    InMux I__2397 (
            .O(N__17103),
            .I(N__17092));
    InMux I__2396 (
            .O(N__17102),
            .I(N__17089));
    InMux I__2395 (
            .O(N__17101),
            .I(N__17086));
    Span4Mux_s2_v I__2394 (
            .O(N__17098),
            .I(N__17081));
    Span4Mux_h I__2393 (
            .O(N__17095),
            .I(N__17081));
    LocalMux I__2392 (
            .O(N__17092),
            .I(N__17078));
    LocalMux I__2391 (
            .O(N__17089),
            .I(\GENERIC_FIFO_1.write_pointer_6 ));
    LocalMux I__2390 (
            .O(N__17086),
            .I(\GENERIC_FIFO_1.write_pointer_6 ));
    Odrv4 I__2389 (
            .O(N__17081),
            .I(\GENERIC_FIFO_1.write_pointer_6 ));
    Odrv12 I__2388 (
            .O(N__17078),
            .I(\GENERIC_FIFO_1.write_pointer_6 ));
    InMux I__2387 (
            .O(N__17069),
            .I(N__17066));
    LocalMux I__2386 (
            .O(N__17066),
            .I(N__17061));
    InMux I__2385 (
            .O(N__17065),
            .I(N__17058));
    InMux I__2384 (
            .O(N__17064),
            .I(N__17053));
    Span4Mux_v I__2383 (
            .O(N__17061),
            .I(N__17047));
    LocalMux I__2382 (
            .O(N__17058),
            .I(N__17047));
    InMux I__2381 (
            .O(N__17057),
            .I(N__17044));
    InMux I__2380 (
            .O(N__17056),
            .I(N__17041));
    LocalMux I__2379 (
            .O(N__17053),
            .I(N__17038));
    InMux I__2378 (
            .O(N__17052),
            .I(N__17035));
    Span4Mux_v I__2377 (
            .O(N__17047),
            .I(N__17030));
    LocalMux I__2376 (
            .O(N__17044),
            .I(N__17030));
    LocalMux I__2375 (
            .O(N__17041),
            .I(N__17025));
    Span12Mux_s2_v I__2374 (
            .O(N__17038),
            .I(N__17025));
    LocalMux I__2373 (
            .O(N__17035),
            .I(\GENERIC_FIFO_1.read_pointer_0 ));
    Odrv4 I__2372 (
            .O(N__17030),
            .I(\GENERIC_FIFO_1.read_pointer_0 ));
    Odrv12 I__2371 (
            .O(N__17025),
            .I(\GENERIC_FIFO_1.read_pointer_0 ));
    CascadeMux I__2370 (
            .O(N__17018),
            .I(N__17015));
    InMux I__2369 (
            .O(N__17015),
            .I(N__17012));
    LocalMux I__2368 (
            .O(N__17012),
            .I(\GENERIC_FIFO_1.n2 ));
    InMux I__2367 (
            .O(N__17009),
            .I(bfn_4_15_0_));
    CascadeMux I__2366 (
            .O(N__17006),
            .I(N__17003));
    InMux I__2365 (
            .O(N__17003),
            .I(N__17000));
    LocalMux I__2364 (
            .O(N__17000),
            .I(\GENERIC_FIFO_1.n1379 ));
    InMux I__2363 (
            .O(N__16997),
            .I(\GENERIC_FIFO_1.n7938 ));
    InMux I__2362 (
            .O(N__16994),
            .I(N__16991));
    LocalMux I__2361 (
            .O(N__16991),
            .I(\GENERIC_FIFO_1.n1391 ));
    CascadeMux I__2360 (
            .O(N__16988),
            .I(N__16985));
    InMux I__2359 (
            .O(N__16985),
            .I(N__16982));
    LocalMux I__2358 (
            .O(N__16982),
            .I(N__16979));
    Odrv12 I__2357 (
            .O(N__16979),
            .I(\GENERIC_FIFO_1.n1378 ));
    InMux I__2356 (
            .O(N__16976),
            .I(N__16973));
    LocalMux I__2355 (
            .O(N__16973),
            .I(N__16970));
    Span4Mux_s3_h I__2354 (
            .O(N__16970),
            .I(N__16967));
    Span4Mux_v I__2353 (
            .O(N__16967),
            .I(N__16964));
    Odrv4 I__2352 (
            .O(N__16964),
            .I(\GENERIC_FIFO_1.n8634 ));
    InMux I__2351 (
            .O(N__16961),
            .I(\GENERIC_FIFO_1.n7939 ));
    CascadeMux I__2350 (
            .O(N__16958),
            .I(N__16955));
    InMux I__2349 (
            .O(N__16955),
            .I(N__16952));
    LocalMux I__2348 (
            .O(N__16952),
            .I(\GENERIC_FIFO_1.n1377 ));
    InMux I__2347 (
            .O(N__16949),
            .I(\GENERIC_FIFO_1.n7940 ));
    InMux I__2346 (
            .O(N__16946),
            .I(N__16943));
    LocalMux I__2345 (
            .O(N__16943),
            .I(\GENERIC_FIFO_1.n1390 ));
    CascadeMux I__2344 (
            .O(N__16940),
            .I(N__16937));
    InMux I__2343 (
            .O(N__16937),
            .I(N__16934));
    LocalMux I__2342 (
            .O(N__16934),
            .I(N__16931));
    Span4Mux_v I__2341 (
            .O(N__16931),
            .I(N__16928));
    Odrv4 I__2340 (
            .O(N__16928),
            .I(\GENERIC_FIFO_1.n1376 ));
    InMux I__2339 (
            .O(N__16925),
            .I(N__16922));
    LocalMux I__2338 (
            .O(N__16922),
            .I(N__16919));
    Span4Mux_s3_h I__2337 (
            .O(N__16919),
            .I(N__16916));
    Span4Mux_v I__2336 (
            .O(N__16916),
            .I(N__16913));
    Odrv4 I__2335 (
            .O(N__16913),
            .I(\GENERIC_FIFO_1.n8628 ));
    InMux I__2334 (
            .O(N__16910),
            .I(\GENERIC_FIFO_1.n7941 ));
    InMux I__2333 (
            .O(N__16907),
            .I(N__16904));
    LocalMux I__2332 (
            .O(N__16904),
            .I(N__16901));
    Span4Mux_s2_v I__2331 (
            .O(N__16901),
            .I(N__16898));
    Odrv4 I__2330 (
            .O(N__16898),
            .I(\GENERIC_FIFO_1.n1375 ));
    InMux I__2329 (
            .O(N__16895),
            .I(\GENERIC_FIFO_1.n7942 ));
    InMux I__2328 (
            .O(N__16892),
            .I(N__16889));
    LocalMux I__2327 (
            .O(N__16889),
            .I(\GENERIC_FIFO_1.n1386 ));
    CascadeMux I__2326 (
            .O(N__16886),
            .I(N__16883));
    InMux I__2325 (
            .O(N__16883),
            .I(N__16880));
    LocalMux I__2324 (
            .O(N__16880),
            .I(\GENERIC_FIFO_1.n1374 ));
    InMux I__2323 (
            .O(N__16877),
            .I(N__16874));
    LocalMux I__2322 (
            .O(N__16874),
            .I(N__16871));
    Span12Mux_v I__2321 (
            .O(N__16871),
            .I(N__16868));
    Odrv12 I__2320 (
            .O(N__16868),
            .I(\GENERIC_FIFO_1.n8632 ));
    InMux I__2319 (
            .O(N__16865),
            .I(\GENERIC_FIFO_1.n7943 ));
    CascadeMux I__2318 (
            .O(N__16862),
            .I(N__16859));
    InMux I__2317 (
            .O(N__16859),
            .I(N__16856));
    LocalMux I__2316 (
            .O(N__16856),
            .I(N__16853));
    Span4Mux_s3_h I__2315 (
            .O(N__16853),
            .I(N__16850));
    Odrv4 I__2314 (
            .O(N__16850),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_7 ));
    InMux I__2313 (
            .O(N__16847),
            .I(N__16844));
    LocalMux I__2312 (
            .O(N__16844),
            .I(\GENERIC_FIFO_1.n17_adj_1280 ));
    InMux I__2311 (
            .O(N__16841),
            .I(N__16838));
    LocalMux I__2310 (
            .O(N__16838),
            .I(N__16835));
    Odrv4 I__2309 (
            .O(N__16835),
            .I(\GENERIC_FIFO_1.n1421 ));
    InMux I__2308 (
            .O(N__16832),
            .I(N__16829));
    LocalMux I__2307 (
            .O(N__16829),
            .I(N__16826));
    Odrv4 I__2306 (
            .O(N__16826),
            .I(\GENERIC_FIFO_1.n1423 ));
    InMux I__2305 (
            .O(N__16823),
            .I(N__16819));
    SRMux I__2304 (
            .O(N__16822),
            .I(N__16816));
    LocalMux I__2303 (
            .O(N__16819),
            .I(N__16808));
    LocalMux I__2302 (
            .O(N__16816),
            .I(N__16808));
    SRMux I__2301 (
            .O(N__16815),
            .I(N__16805));
    SRMux I__2300 (
            .O(N__16814),
            .I(N__16799));
    InMux I__2299 (
            .O(N__16813),
            .I(N__16796));
    Span4Mux_s3_v I__2298 (
            .O(N__16808),
            .I(N__16784));
    LocalMux I__2297 (
            .O(N__16805),
            .I(N__16784));
    CascadeMux I__2296 (
            .O(N__16804),
            .I(N__16780));
    InMux I__2295 (
            .O(N__16803),
            .I(N__16773));
    InMux I__2294 (
            .O(N__16802),
            .I(N__16773));
    LocalMux I__2293 (
            .O(N__16799),
            .I(N__16770));
    LocalMux I__2292 (
            .O(N__16796),
            .I(N__16767));
    InMux I__2291 (
            .O(N__16795),
            .I(N__16752));
    InMux I__2290 (
            .O(N__16794),
            .I(N__16752));
    InMux I__2289 (
            .O(N__16793),
            .I(N__16752));
    InMux I__2288 (
            .O(N__16792),
            .I(N__16752));
    InMux I__2287 (
            .O(N__16791),
            .I(N__16752));
    InMux I__2286 (
            .O(N__16790),
            .I(N__16752));
    InMux I__2285 (
            .O(N__16789),
            .I(N__16752));
    Span4Mux_v I__2284 (
            .O(N__16784),
            .I(N__16749));
    InMux I__2283 (
            .O(N__16783),
            .I(N__16740));
    InMux I__2282 (
            .O(N__16780),
            .I(N__16740));
    InMux I__2281 (
            .O(N__16779),
            .I(N__16740));
    InMux I__2280 (
            .O(N__16778),
            .I(N__16740));
    LocalMux I__2279 (
            .O(N__16773),
            .I(N__16737));
    Sp12to4 I__2278 (
            .O(N__16770),
            .I(N__16732));
    Span12Mux_s11_h I__2277 (
            .O(N__16767),
            .I(N__16732));
    LocalMux I__2276 (
            .O(N__16752),
            .I(writeByte));
    Odrv4 I__2275 (
            .O(N__16749),
            .I(writeByte));
    LocalMux I__2274 (
            .O(N__16740),
            .I(writeByte));
    Odrv4 I__2273 (
            .O(N__16737),
            .I(writeByte));
    Odrv12 I__2272 (
            .O(N__16732),
            .I(writeByte));
    InMux I__2271 (
            .O(N__16721),
            .I(N__16718));
    LocalMux I__2270 (
            .O(N__16718),
            .I(N__16714));
    InMux I__2269 (
            .O(N__16717),
            .I(N__16711));
    Span4Mux_v I__2268 (
            .O(N__16714),
            .I(N__16708));
    LocalMux I__2267 (
            .O(N__16711),
            .I(N__16703));
    Span4Mux_v I__2266 (
            .O(N__16708),
            .I(N__16700));
    InMux I__2265 (
            .O(N__16707),
            .I(N__16695));
    InMux I__2264 (
            .O(N__16706),
            .I(N__16695));
    Odrv4 I__2263 (
            .O(N__16703),
            .I(n9));
    Odrv4 I__2262 (
            .O(N__16700),
            .I(n9));
    LocalMux I__2261 (
            .O(N__16695),
            .I(n9));
    SRMux I__2260 (
            .O(N__16688),
            .I(N__16682));
    SRMux I__2259 (
            .O(N__16687),
            .I(N__16679));
    CEMux I__2258 (
            .O(N__16686),
            .I(N__16676));
    CEMux I__2257 (
            .O(N__16685),
            .I(N__16673));
    LocalMux I__2256 (
            .O(N__16682),
            .I(N__16670));
    LocalMux I__2255 (
            .O(N__16679),
            .I(N__16667));
    LocalMux I__2254 (
            .O(N__16676),
            .I(N__16664));
    LocalMux I__2253 (
            .O(N__16673),
            .I(N__16661));
    Span4Mux_s3_h I__2252 (
            .O(N__16670),
            .I(N__16658));
    Span4Mux_s3_h I__2251 (
            .O(N__16667),
            .I(N__16655));
    Span12Mux_s3_h I__2250 (
            .O(N__16664),
            .I(N__16652));
    Span4Mux_h I__2249 (
            .O(N__16661),
            .I(N__16649));
    Span4Mux_v I__2248 (
            .O(N__16658),
            .I(N__16646));
    Span4Mux_v I__2247 (
            .O(N__16655),
            .I(N__16643));
    Odrv12 I__2246 (
            .O(N__16652),
            .I(\Inst_eia232.Inst_transmitter.n3608 ));
    Odrv4 I__2245 (
            .O(N__16649),
            .I(\Inst_eia232.Inst_transmitter.n3608 ));
    Odrv4 I__2244 (
            .O(N__16646),
            .I(\Inst_eia232.Inst_transmitter.n3608 ));
    Odrv4 I__2243 (
            .O(N__16643),
            .I(\Inst_eia232.Inst_transmitter.n3608 ));
    CascadeMux I__2242 (
            .O(N__16634),
            .I(N__16631));
    CascadeBuf I__2241 (
            .O(N__16631),
            .I(N__16626));
    CascadeMux I__2240 (
            .O(N__16630),
            .I(N__16623));
    InMux I__2239 (
            .O(N__16629),
            .I(N__16620));
    CascadeMux I__2238 (
            .O(N__16626),
            .I(N__16617));
    InMux I__2237 (
            .O(N__16623),
            .I(N__16612));
    LocalMux I__2236 (
            .O(N__16620),
            .I(N__16609));
    InMux I__2235 (
            .O(N__16617),
            .I(N__16606));
    InMux I__2234 (
            .O(N__16616),
            .I(N__16603));
    InMux I__2233 (
            .O(N__16615),
            .I(N__16600));
    LocalMux I__2232 (
            .O(N__16612),
            .I(N__16597));
    Span4Mux_v I__2231 (
            .O(N__16609),
            .I(N__16592));
    LocalMux I__2230 (
            .O(N__16606),
            .I(N__16592));
    LocalMux I__2229 (
            .O(N__16603),
            .I(\GENERIC_FIFO_1.write_pointer_0 ));
    LocalMux I__2228 (
            .O(N__16600),
            .I(\GENERIC_FIFO_1.write_pointer_0 ));
    Odrv12 I__2227 (
            .O(N__16597),
            .I(\GENERIC_FIFO_1.write_pointer_0 ));
    Odrv4 I__2226 (
            .O(N__16592),
            .I(\GENERIC_FIFO_1.write_pointer_0 ));
    CascadeMux I__2225 (
            .O(N__16583),
            .I(N__16580));
    CascadeBuf I__2224 (
            .O(N__16580),
            .I(N__16576));
    InMux I__2223 (
            .O(N__16579),
            .I(N__16572));
    CascadeMux I__2222 (
            .O(N__16576),
            .I(N__16569));
    InMux I__2221 (
            .O(N__16575),
            .I(N__16564));
    LocalMux I__2220 (
            .O(N__16572),
            .I(N__16561));
    InMux I__2219 (
            .O(N__16569),
            .I(N__16558));
    InMux I__2218 (
            .O(N__16568),
            .I(N__16555));
    InMux I__2217 (
            .O(N__16567),
            .I(N__16552));
    LocalMux I__2216 (
            .O(N__16564),
            .I(N__16549));
    Span4Mux_v I__2215 (
            .O(N__16561),
            .I(N__16544));
    LocalMux I__2214 (
            .O(N__16558),
            .I(N__16544));
    LocalMux I__2213 (
            .O(N__16555),
            .I(\GENERIC_FIFO_1.write_pointer_1 ));
    LocalMux I__2212 (
            .O(N__16552),
            .I(\GENERIC_FIFO_1.write_pointer_1 ));
    Odrv12 I__2211 (
            .O(N__16549),
            .I(\GENERIC_FIFO_1.write_pointer_1 ));
    Odrv4 I__2210 (
            .O(N__16544),
            .I(\GENERIC_FIFO_1.write_pointer_1 ));
    CascadeMux I__2209 (
            .O(N__16535),
            .I(N__16532));
    CascadeBuf I__2208 (
            .O(N__16532),
            .I(N__16527));
    InMux I__2207 (
            .O(N__16531),
            .I(N__16524));
    InMux I__2206 (
            .O(N__16530),
            .I(N__16521));
    CascadeMux I__2205 (
            .O(N__16527),
            .I(N__16518));
    LocalMux I__2204 (
            .O(N__16524),
            .I(N__16513));
    LocalMux I__2203 (
            .O(N__16521),
            .I(N__16510));
    InMux I__2202 (
            .O(N__16518),
            .I(N__16507));
    InMux I__2201 (
            .O(N__16517),
            .I(N__16504));
    InMux I__2200 (
            .O(N__16516),
            .I(N__16501));
    Span4Mux_v I__2199 (
            .O(N__16513),
            .I(N__16494));
    Span4Mux_v I__2198 (
            .O(N__16510),
            .I(N__16494));
    LocalMux I__2197 (
            .O(N__16507),
            .I(N__16494));
    LocalMux I__2196 (
            .O(N__16504),
            .I(\GENERIC_FIFO_1.write_pointer_2 ));
    LocalMux I__2195 (
            .O(N__16501),
            .I(\GENERIC_FIFO_1.write_pointer_2 ));
    Odrv4 I__2194 (
            .O(N__16494),
            .I(\GENERIC_FIFO_1.write_pointer_2 ));
    CascadeMux I__2193 (
            .O(N__16487),
            .I(N__16484));
    CascadeBuf I__2192 (
            .O(N__16484),
            .I(N__16479));
    InMux I__2191 (
            .O(N__16483),
            .I(N__16476));
    InMux I__2190 (
            .O(N__16482),
            .I(N__16473));
    CascadeMux I__2189 (
            .O(N__16479),
            .I(N__16470));
    LocalMux I__2188 (
            .O(N__16476),
            .I(N__16465));
    LocalMux I__2187 (
            .O(N__16473),
            .I(N__16462));
    InMux I__2186 (
            .O(N__16470),
            .I(N__16459));
    InMux I__2185 (
            .O(N__16469),
            .I(N__16456));
    InMux I__2184 (
            .O(N__16468),
            .I(N__16453));
    Span4Mux_v I__2183 (
            .O(N__16465),
            .I(N__16446));
    Span4Mux_v I__2182 (
            .O(N__16462),
            .I(N__16446));
    LocalMux I__2181 (
            .O(N__16459),
            .I(N__16446));
    LocalMux I__2180 (
            .O(N__16456),
            .I(\GENERIC_FIFO_1.write_pointer_3 ));
    LocalMux I__2179 (
            .O(N__16453),
            .I(\GENERIC_FIFO_1.write_pointer_3 ));
    Odrv4 I__2178 (
            .O(N__16446),
            .I(\GENERIC_FIFO_1.write_pointer_3 ));
    CascadeMux I__2177 (
            .O(N__16439),
            .I(N__16436));
    CascadeBuf I__2176 (
            .O(N__16436),
            .I(N__16433));
    CascadeMux I__2175 (
            .O(N__16433),
            .I(N__16430));
    InMux I__2174 (
            .O(N__16430),
            .I(N__16427));
    LocalMux I__2173 (
            .O(N__16427),
            .I(\GENERIC_FIFO_1.n76 ));
    CascadeMux I__2172 (
            .O(N__16424),
            .I(N__16421));
    CascadeBuf I__2171 (
            .O(N__16421),
            .I(N__16418));
    CascadeMux I__2170 (
            .O(N__16418),
            .I(N__16415));
    InMux I__2169 (
            .O(N__16415),
            .I(N__16412));
    LocalMux I__2168 (
            .O(N__16412),
            .I(\GENERIC_FIFO_1.n75 ));
    CascadeMux I__2167 (
            .O(N__16409),
            .I(N__16406));
    CascadeBuf I__2166 (
            .O(N__16406),
            .I(N__16403));
    CascadeMux I__2165 (
            .O(N__16403),
            .I(N__16400));
    InMux I__2164 (
            .O(N__16400),
            .I(N__16397));
    LocalMux I__2163 (
            .O(N__16397),
            .I(\GENERIC_FIFO_1.n74 ));
    CascadeMux I__2162 (
            .O(N__16394),
            .I(N__16391));
    CascadeBuf I__2161 (
            .O(N__16391),
            .I(N__16388));
    CascadeMux I__2160 (
            .O(N__16388),
            .I(N__16385));
    InMux I__2159 (
            .O(N__16385),
            .I(N__16382));
    LocalMux I__2158 (
            .O(N__16382),
            .I(\GENERIC_FIFO_1.n73 ));
    InMux I__2157 (
            .O(N__16379),
            .I(N__16376));
    LocalMux I__2156 (
            .O(N__16376),
            .I(N__16373));
    Span4Mux_v I__2155 (
            .O(N__16373),
            .I(N__16370));
    Odrv4 I__2154 (
            .O(N__16370),
            .I(\GENERIC_FIFO_1.n1420 ));
    CascadeMux I__2153 (
            .O(N__16367),
            .I(N__16364));
    CascadeBuf I__2152 (
            .O(N__16364),
            .I(N__16361));
    CascadeMux I__2151 (
            .O(N__16361),
            .I(N__16358));
    InMux I__2150 (
            .O(N__16358),
            .I(N__16355));
    LocalMux I__2149 (
            .O(N__16355),
            .I(\GENERIC_FIFO_1.n72 ));
    CascadeMux I__2148 (
            .O(N__16352),
            .I(\GENERIC_FIFO_1.n16_adj_1279_cascade_ ));
    InMux I__2147 (
            .O(N__16349),
            .I(N__16331));
    InMux I__2146 (
            .O(N__16348),
            .I(N__16331));
    InMux I__2145 (
            .O(N__16347),
            .I(N__16331));
    InMux I__2144 (
            .O(N__16346),
            .I(N__16331));
    InMux I__2143 (
            .O(N__16345),
            .I(N__16328));
    InMux I__2142 (
            .O(N__16344),
            .I(N__16325));
    InMux I__2141 (
            .O(N__16343),
            .I(N__16316));
    InMux I__2140 (
            .O(N__16342),
            .I(N__16316));
    InMux I__2139 (
            .O(N__16341),
            .I(N__16316));
    InMux I__2138 (
            .O(N__16340),
            .I(N__16316));
    LocalMux I__2137 (
            .O(N__16331),
            .I(N__16313));
    LocalMux I__2136 (
            .O(N__16328),
            .I(N__16308));
    LocalMux I__2135 (
            .O(N__16325),
            .I(N__16308));
    LocalMux I__2134 (
            .O(N__16316),
            .I(N__16305));
    Span4Mux_v I__2133 (
            .O(N__16313),
            .I(N__16302));
    Span4Mux_s2_h I__2132 (
            .O(N__16308),
            .I(N__16297));
    Span4Mux_v I__2131 (
            .O(N__16305),
            .I(N__16297));
    Span4Mux_v I__2130 (
            .O(N__16302),
            .I(N__16292));
    Span4Mux_v I__2129 (
            .O(N__16297),
            .I(N__16292));
    Odrv4 I__2128 (
            .O(N__16292),
            .I(\GENERIC_FIFO_1.n142 ));
    CascadeMux I__2127 (
            .O(N__16289),
            .I(N__16286));
    InMux I__2126 (
            .O(N__16286),
            .I(N__16283));
    LocalMux I__2125 (
            .O(N__16283),
            .I(N__16280));
    Span4Mux_v I__2124 (
            .O(N__16280),
            .I(N__16277));
    Odrv4 I__2123 (
            .O(N__16277),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_7 ));
    SRMux I__2122 (
            .O(N__16274),
            .I(N__16271));
    LocalMux I__2121 (
            .O(N__16271),
            .I(N__16268));
    Span4Mux_s2_v I__2120 (
            .O(N__16268),
            .I(N__16265));
    Span4Mux_v I__2119 (
            .O(N__16265),
            .I(N__16262));
    Odrv4 I__2118 (
            .O(N__16262),
            .I(\Inst_eia232.Inst_receiver.n4628 ));
    InMux I__2117 (
            .O(N__16259),
            .I(N__16256));
    LocalMux I__2116 (
            .O(N__16256),
            .I(N__16253));
    Span4Mux_v I__2115 (
            .O(N__16253),
            .I(N__16250));
    Span4Mux_h I__2114 (
            .O(N__16250),
            .I(N__16246));
    InMux I__2113 (
            .O(N__16249),
            .I(N__16243));
    Span4Mux_v I__2112 (
            .O(N__16246),
            .I(N__16238));
    LocalMux I__2111 (
            .O(N__16243),
            .I(N__16238));
    Span4Mux_v I__2110 (
            .O(N__16238),
            .I(N__16235));
    Odrv4 I__2109 (
            .O(N__16235),
            .I(\Inst_eia232.Inst_transmitter.paused ));
    SRMux I__2108 (
            .O(N__16232),
            .I(N__16229));
    LocalMux I__2107 (
            .O(N__16229),
            .I(N__16225));
    SRMux I__2106 (
            .O(N__16228),
            .I(N__16222));
    Span4Mux_s2_h I__2105 (
            .O(N__16225),
            .I(N__16217));
    LocalMux I__2104 (
            .O(N__16222),
            .I(N__16217));
    Span4Mux_v I__2103 (
            .O(N__16217),
            .I(N__16214));
    Span4Mux_v I__2102 (
            .O(N__16214),
            .I(N__16211));
    Odrv4 I__2101 (
            .O(N__16211),
            .I(\Inst_eia232.Inst_transmitter.n4634 ));
    SRMux I__2100 (
            .O(N__16208),
            .I(N__16199));
    InMux I__2099 (
            .O(N__16207),
            .I(N__16199));
    InMux I__2098 (
            .O(N__16206),
            .I(N__16199));
    LocalMux I__2097 (
            .O(N__16199),
            .I(N__16193));
    CascadeMux I__2096 (
            .O(N__16198),
            .I(N__16188));
    InMux I__2095 (
            .O(N__16197),
            .I(N__16182));
    InMux I__2094 (
            .O(N__16196),
            .I(N__16182));
    Span4Mux_h I__2093 (
            .O(N__16193),
            .I(N__16179));
    InMux I__2092 (
            .O(N__16192),
            .I(N__16174));
    InMux I__2091 (
            .O(N__16191),
            .I(N__16170));
    InMux I__2090 (
            .O(N__16188),
            .I(N__16165));
    InMux I__2089 (
            .O(N__16187),
            .I(N__16165));
    LocalMux I__2088 (
            .O(N__16182),
            .I(N__16160));
    Span4Mux_v I__2087 (
            .O(N__16179),
            .I(N__16160));
    InMux I__2086 (
            .O(N__16178),
            .I(N__16155));
    InMux I__2085 (
            .O(N__16177),
            .I(N__16155));
    LocalMux I__2084 (
            .O(N__16174),
            .I(N__16152));
    InMux I__2083 (
            .O(N__16173),
            .I(N__16149));
    LocalMux I__2082 (
            .O(N__16170),
            .I(state_0));
    LocalMux I__2081 (
            .O(N__16165),
            .I(state_0));
    Odrv4 I__2080 (
            .O(N__16160),
            .I(state_0));
    LocalMux I__2079 (
            .O(N__16155),
            .I(state_0));
    Odrv4 I__2078 (
            .O(N__16152),
            .I(state_0));
    LocalMux I__2077 (
            .O(N__16149),
            .I(state_0));
    InMux I__2076 (
            .O(N__16136),
            .I(N__16133));
    LocalMux I__2075 (
            .O(N__16133),
            .I(N__16125));
    CascadeMux I__2074 (
            .O(N__16132),
            .I(N__16122));
    InMux I__2073 (
            .O(N__16131),
            .I(N__16112));
    InMux I__2072 (
            .O(N__16130),
            .I(N__16112));
    InMux I__2071 (
            .O(N__16129),
            .I(N__16112));
    InMux I__2070 (
            .O(N__16128),
            .I(N__16112));
    Span4Mux_h I__2069 (
            .O(N__16125),
            .I(N__16109));
    InMux I__2068 (
            .O(N__16122),
            .I(N__16104));
    InMux I__2067 (
            .O(N__16121),
            .I(N__16104));
    LocalMux I__2066 (
            .O(N__16112),
            .I(N__16101));
    Span4Mux_v I__2065 (
            .O(N__16109),
            .I(N__16098));
    LocalMux I__2064 (
            .O(N__16104),
            .I(\Inst_eia232.Inst_transmitter.n2580 ));
    Odrv4 I__2063 (
            .O(N__16101),
            .I(\Inst_eia232.Inst_transmitter.n2580 ));
    Odrv4 I__2062 (
            .O(N__16098),
            .I(\Inst_eia232.Inst_transmitter.n2580 ));
    InMux I__2061 (
            .O(N__16091),
            .I(N__16088));
    LocalMux I__2060 (
            .O(N__16088),
            .I(N__16084));
    InMux I__2059 (
            .O(N__16087),
            .I(N__16081));
    Span4Mux_s2_h I__2058 (
            .O(N__16084),
            .I(N__16076));
    LocalMux I__2057 (
            .O(N__16081),
            .I(N__16076));
    Span4Mux_v I__2056 (
            .O(N__16076),
            .I(N__16073));
    Odrv4 I__2055 (
            .O(N__16073),
            .I(\Inst_eia232.Inst_transmitter.n8527 ));
    CascadeMux I__2054 (
            .O(N__16070),
            .I(N__16065));
    CascadeMux I__2053 (
            .O(N__16069),
            .I(N__16062));
    InMux I__2052 (
            .O(N__16068),
            .I(N__16059));
    InMux I__2051 (
            .O(N__16065),
            .I(N__16056));
    InMux I__2050 (
            .O(N__16062),
            .I(N__16053));
    LocalMux I__2049 (
            .O(N__16059),
            .I(N__16050));
    LocalMux I__2048 (
            .O(N__16056),
            .I(N__16047));
    LocalMux I__2047 (
            .O(N__16053),
            .I(N__16044));
    Span4Mux_v I__2046 (
            .O(N__16050),
            .I(N__16039));
    Span4Mux_s3_h I__2045 (
            .O(N__16047),
            .I(N__16039));
    Span4Mux_h I__2044 (
            .O(N__16044),
            .I(N__16036));
    Odrv4 I__2043 (
            .O(N__16039),
            .I(\Inst_eia232.id ));
    Odrv4 I__2042 (
            .O(N__16036),
            .I(\Inst_eia232.id ));
    InMux I__2041 (
            .O(N__16031),
            .I(N__16028));
    LocalMux I__2040 (
            .O(N__16028),
            .I(N__16025));
    Span4Mux_v I__2039 (
            .O(N__16025),
            .I(N__16022));
    Span4Mux_v I__2038 (
            .O(N__16022),
            .I(N__16019));
    Odrv4 I__2037 (
            .O(N__16019),
            .I(\Inst_eia232.Inst_transmitter.n971 ));
    InMux I__2036 (
            .O(N__16016),
            .I(N__16007));
    InMux I__2035 (
            .O(N__16015),
            .I(N__16007));
    InMux I__2034 (
            .O(N__16014),
            .I(N__16000));
    InMux I__2033 (
            .O(N__16013),
            .I(N__16000));
    InMux I__2032 (
            .O(N__16012),
            .I(N__16000));
    LocalMux I__2031 (
            .O(N__16007),
            .I(N__15992));
    LocalMux I__2030 (
            .O(N__16000),
            .I(N__15992));
    InMux I__2029 (
            .O(N__15999),
            .I(N__15977));
    InMux I__2028 (
            .O(N__15998),
            .I(N__15974));
    InMux I__2027 (
            .O(N__15997),
            .I(N__15971));
    Span4Mux_v I__2026 (
            .O(N__15992),
            .I(N__15968));
    InMux I__2025 (
            .O(N__15991),
            .I(N__15952));
    InMux I__2024 (
            .O(N__15990),
            .I(N__15952));
    InMux I__2023 (
            .O(N__15989),
            .I(N__15952));
    InMux I__2022 (
            .O(N__15988),
            .I(N__15952));
    InMux I__2021 (
            .O(N__15987),
            .I(N__15952));
    InMux I__2020 (
            .O(N__15986),
            .I(N__15952));
    InMux I__2019 (
            .O(N__15985),
            .I(N__15952));
    InMux I__2018 (
            .O(N__15984),
            .I(N__15948));
    InMux I__2017 (
            .O(N__15983),
            .I(N__15939));
    InMux I__2016 (
            .O(N__15982),
            .I(N__15939));
    InMux I__2015 (
            .O(N__15981),
            .I(N__15939));
    InMux I__2014 (
            .O(N__15980),
            .I(N__15939));
    LocalMux I__2013 (
            .O(N__15977),
            .I(N__15936));
    LocalMux I__2012 (
            .O(N__15974),
            .I(N__15931));
    LocalMux I__2011 (
            .O(N__15971),
            .I(N__15931));
    Span4Mux_v I__2010 (
            .O(N__15968),
            .I(N__15928));
    InMux I__2009 (
            .O(N__15967),
            .I(N__15925));
    LocalMux I__2008 (
            .O(N__15952),
            .I(N__15922));
    InMux I__2007 (
            .O(N__15951),
            .I(N__15919));
    LocalMux I__2006 (
            .O(N__15948),
            .I(state_1));
    LocalMux I__2005 (
            .O(N__15939),
            .I(state_1));
    Odrv4 I__2004 (
            .O(N__15936),
            .I(state_1));
    Odrv12 I__2003 (
            .O(N__15931),
            .I(state_1));
    Odrv4 I__2002 (
            .O(N__15928),
            .I(state_1));
    LocalMux I__2001 (
            .O(N__15925),
            .I(state_1));
    Odrv4 I__2000 (
            .O(N__15922),
            .I(state_1));
    LocalMux I__1999 (
            .O(N__15919),
            .I(state_1));
    SRMux I__1998 (
            .O(N__15902),
            .I(N__15899));
    LocalMux I__1997 (
            .O(N__15899),
            .I(N__15896));
    Span4Mux_v I__1996 (
            .O(N__15896),
            .I(N__15893));
    Span4Mux_s0_h I__1995 (
            .O(N__15893),
            .I(N__15890));
    Odrv4 I__1994 (
            .O(N__15890),
            .I(\Inst_eia232.Inst_transmitter.n4712 ));
    CascadeMux I__1993 (
            .O(N__15887),
            .I(N__15884));
    CascadeBuf I__1992 (
            .O(N__15884),
            .I(N__15881));
    CascadeMux I__1991 (
            .O(N__15881),
            .I(N__15878));
    InMux I__1990 (
            .O(N__15878),
            .I(N__15875));
    LocalMux I__1989 (
            .O(N__15875),
            .I(\GENERIC_FIFO_1.n77 ));
    InMux I__1988 (
            .O(N__15872),
            .I(N__15868));
    CascadeMux I__1987 (
            .O(N__15871),
            .I(N__15865));
    LocalMux I__1986 (
            .O(N__15868),
            .I(N__15861));
    InMux I__1985 (
            .O(N__15865),
            .I(N__15856));
    InMux I__1984 (
            .O(N__15864),
            .I(N__15856));
    Odrv4 I__1983 (
            .O(N__15861),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0 ));
    LocalMux I__1982 (
            .O(N__15856),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0 ));
    InMux I__1981 (
            .O(N__15851),
            .I(N__15848));
    LocalMux I__1980 (
            .O(N__15848),
            .I(N__15844));
    CascadeMux I__1979 (
            .O(N__15847),
            .I(N__15841));
    Span4Mux_v I__1978 (
            .O(N__15844),
            .I(N__15837));
    InMux I__1977 (
            .O(N__15841),
            .I(N__15832));
    InMux I__1976 (
            .O(N__15840),
            .I(N__15832));
    Odrv4 I__1975 (
            .O(N__15837),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4 ));
    LocalMux I__1974 (
            .O(N__15832),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4 ));
    InMux I__1973 (
            .O(N__15827),
            .I(N__15824));
    LocalMux I__1972 (
            .O(N__15824),
            .I(N__15821));
    Span4Mux_v I__1971 (
            .O(N__15821),
            .I(N__15818));
    Span4Mux_s1_h I__1970 (
            .O(N__15818),
            .I(N__15813));
    InMux I__1969 (
            .O(N__15817),
            .I(N__15808));
    InMux I__1968 (
            .O(N__15816),
            .I(N__15808));
    Odrv4 I__1967 (
            .O(N__15813),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5 ));
    LocalMux I__1966 (
            .O(N__15808),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5 ));
    CascadeMux I__1965 (
            .O(N__15803),
            .I(N__15800));
    InMux I__1964 (
            .O(N__15800),
            .I(N__15797));
    LocalMux I__1963 (
            .O(N__15797),
            .I(N__15794));
    Span12Mux_s7_v I__1962 (
            .O(N__15794),
            .I(N__15790));
    InMux I__1961 (
            .O(N__15793),
            .I(N__15787));
    Odrv12 I__1960 (
            .O(N__15790),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6 ));
    LocalMux I__1959 (
            .O(N__15787),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6 ));
    CascadeMux I__1958 (
            .O(N__15782),
            .I(N__15779));
    CascadeBuf I__1957 (
            .O(N__15779),
            .I(N__15776));
    CascadeMux I__1956 (
            .O(N__15776),
            .I(N__15773));
    InMux I__1955 (
            .O(N__15773),
            .I(N__15770));
    LocalMux I__1954 (
            .O(N__15770),
            .I(N__15767));
    Span4Mux_s3_h I__1953 (
            .O(N__15767),
            .I(N__15764));
    Odrv4 I__1952 (
            .O(N__15764),
            .I(\GENERIC_FIFO_1.n71 ));
    CascadeMux I__1951 (
            .O(N__15761),
            .I(N__15758));
    CascadeBuf I__1950 (
            .O(N__15758),
            .I(N__15755));
    CascadeMux I__1949 (
            .O(N__15755),
            .I(N__15752));
    InMux I__1948 (
            .O(N__15752),
            .I(N__15749));
    LocalMux I__1947 (
            .O(N__15749),
            .I(N__15746));
    Span4Mux_v I__1946 (
            .O(N__15746),
            .I(N__15743));
    Odrv4 I__1945 (
            .O(N__15743),
            .I(\GENERIC_FIFO_1.n70 ));
    InMux I__1944 (
            .O(N__15740),
            .I(N__15737));
    LocalMux I__1943 (
            .O(N__15737),
            .I(N__15733));
    InMux I__1942 (
            .O(N__15736),
            .I(N__15730));
    Span4Mux_v I__1941 (
            .O(N__15733),
            .I(N__15727));
    LocalMux I__1940 (
            .O(N__15730),
            .I(N__15724));
    Odrv4 I__1939 (
            .O(N__15727),
            .I(\GENERIC_FIFO_1.n8779 ));
    Odrv12 I__1938 (
            .O(N__15724),
            .I(\GENERIC_FIFO_1.n8779 ));
    InMux I__1937 (
            .O(N__15719),
            .I(N__15715));
    InMux I__1936 (
            .O(N__15718),
            .I(N__15712));
    LocalMux I__1935 (
            .O(N__15715),
            .I(valueRegister_0));
    LocalMux I__1934 (
            .O(N__15712),
            .I(valueRegister_0));
    CascadeMux I__1933 (
            .O(N__15707),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_cascade_ ));
    CascadeMux I__1932 (
            .O(N__15704),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9114_cascade_ ));
    InMux I__1931 (
            .O(N__15701),
            .I(N__15698));
    LocalMux I__1930 (
            .O(N__15698),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_0 ));
    InMux I__1929 (
            .O(N__15695),
            .I(N__15692));
    LocalMux I__1928 (
            .O(N__15692),
            .I(N__15689));
    Span4Mux_s3_h I__1927 (
            .O(N__15689),
            .I(N__15686));
    Odrv4 I__1926 (
            .O(N__15686),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7 ));
    CascadeMux I__1925 (
            .O(N__15683),
            .I(N__15680));
    InMux I__1924 (
            .O(N__15680),
            .I(N__15677));
    LocalMux I__1923 (
            .O(N__15677),
            .I(N__15674));
    Span4Mux_h I__1922 (
            .O(N__15674),
            .I(N__15671));
    Odrv4 I__1921 (
            .O(N__15671),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9108 ));
    InMux I__1920 (
            .O(N__15668),
            .I(N__15664));
    InMux I__1919 (
            .O(N__15667),
            .I(N__15661));
    LocalMux I__1918 (
            .O(N__15664),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16 ));
    LocalMux I__1917 (
            .O(N__15661),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16 ));
    CascadeMux I__1916 (
            .O(N__15656),
            .I(N__15652));
    InMux I__1915 (
            .O(N__15655),
            .I(N__15648));
    InMux I__1914 (
            .O(N__15652),
            .I(N__15645));
    InMux I__1913 (
            .O(N__15651),
            .I(N__15642));
    LocalMux I__1912 (
            .O(N__15648),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16 ));
    LocalMux I__1911 (
            .O(N__15645),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16 ));
    LocalMux I__1910 (
            .O(N__15642),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16 ));
    InMux I__1909 (
            .O(N__15635),
            .I(N__15624));
    InMux I__1908 (
            .O(N__15634),
            .I(N__15624));
    InMux I__1907 (
            .O(N__15633),
            .I(N__15624));
    InMux I__1906 (
            .O(N__15632),
            .I(N__15621));
    InMux I__1905 (
            .O(N__15631),
            .I(N__15618));
    LocalMux I__1904 (
            .O(N__15624),
            .I(N__15613));
    LocalMux I__1903 (
            .O(N__15621),
            .I(N__15613));
    LocalMux I__1902 (
            .O(N__15618),
            .I(\Inst_eia232.Inst_receiver.n14_adj_1265 ));
    Odrv4 I__1901 (
            .O(N__15613),
            .I(\Inst_eia232.Inst_receiver.n14_adj_1265 ));
    InMux I__1900 (
            .O(N__15608),
            .I(N__15593));
    InMux I__1899 (
            .O(N__15607),
            .I(N__15593));
    InMux I__1898 (
            .O(N__15606),
            .I(N__15593));
    InMux I__1897 (
            .O(N__15605),
            .I(N__15593));
    InMux I__1896 (
            .O(N__15604),
            .I(N__15593));
    LocalMux I__1895 (
            .O(N__15593),
            .I(\Inst_eia232.Inst_receiver.n112 ));
    CascadeMux I__1894 (
            .O(N__15590),
            .I(\Inst_eia232.Inst_receiver.n112_cascade_ ));
    InMux I__1893 (
            .O(N__15587),
            .I(N__15583));
    InMux I__1892 (
            .O(N__15586),
            .I(N__15580));
    LocalMux I__1891 (
            .O(N__15583),
            .I(N__15577));
    LocalMux I__1890 (
            .O(N__15580),
            .I(\Inst_eia232.Inst_receiver.n90 ));
    Odrv4 I__1889 (
            .O(N__15577),
            .I(\Inst_eia232.Inst_receiver.n90 ));
    InMux I__1888 (
            .O(N__15572),
            .I(N__15563));
    InMux I__1887 (
            .O(N__15571),
            .I(N__15563));
    InMux I__1886 (
            .O(N__15570),
            .I(N__15563));
    LocalMux I__1885 (
            .O(N__15563),
            .I(N__15559));
    InMux I__1884 (
            .O(N__15562),
            .I(N__15556));
    Odrv4 I__1883 (
            .O(N__15559),
            .I(\Inst_eia232.Inst_receiver.n5498 ));
    LocalMux I__1882 (
            .O(N__15556),
            .I(\Inst_eia232.Inst_receiver.n5498 ));
    InMux I__1881 (
            .O(N__15551),
            .I(N__15546));
    CascadeMux I__1880 (
            .O(N__15550),
            .I(N__15542));
    CascadeMux I__1879 (
            .O(N__15549),
            .I(N__15539));
    LocalMux I__1878 (
            .O(N__15546),
            .I(N__15534));
    InMux I__1877 (
            .O(N__15545),
            .I(N__15523));
    InMux I__1876 (
            .O(N__15542),
            .I(N__15523));
    InMux I__1875 (
            .O(N__15539),
            .I(N__15523));
    InMux I__1874 (
            .O(N__15538),
            .I(N__15523));
    InMux I__1873 (
            .O(N__15537),
            .I(N__15523));
    Odrv4 I__1872 (
            .O(N__15534),
            .I(cmd_6));
    LocalMux I__1871 (
            .O(N__15523),
            .I(cmd_6));
    CascadeMux I__1870 (
            .O(N__15518),
            .I(n5698_cascade_));
    InMux I__1869 (
            .O(N__15515),
            .I(N__15512));
    LocalMux I__1868 (
            .O(N__15512),
            .I(N__15503));
    InMux I__1867 (
            .O(N__15511),
            .I(N__15500));
    InMux I__1866 (
            .O(N__15510),
            .I(N__15489));
    InMux I__1865 (
            .O(N__15509),
            .I(N__15489));
    InMux I__1864 (
            .O(N__15508),
            .I(N__15489));
    InMux I__1863 (
            .O(N__15507),
            .I(N__15489));
    InMux I__1862 (
            .O(N__15506),
            .I(N__15489));
    Odrv4 I__1861 (
            .O(N__15503),
            .I(nstate_2_N_241_0));
    LocalMux I__1860 (
            .O(N__15500),
            .I(nstate_2_N_241_0));
    LocalMux I__1859 (
            .O(N__15489),
            .I(nstate_2_N_241_0));
    InMux I__1858 (
            .O(N__15482),
            .I(N__15479));
    LocalMux I__1857 (
            .O(N__15479),
            .I(N__15476));
    Span4Mux_h I__1856 (
            .O(N__15476),
            .I(N__15472));
    InMux I__1855 (
            .O(N__15475),
            .I(N__15469));
    Odrv4 I__1854 (
            .O(N__15472),
            .I(\Inst_eia232.xon ));
    LocalMux I__1853 (
            .O(N__15469),
            .I(\Inst_eia232.xon ));
    CascadeMux I__1852 (
            .O(N__15464),
            .I(\Inst_eia232.Inst_receiver.n75_cascade_ ));
    InMux I__1851 (
            .O(N__15461),
            .I(N__15458));
    LocalMux I__1850 (
            .O(N__15458),
            .I(\Inst_eia232.Inst_receiver.n5597 ));
    CascadeMux I__1849 (
            .O(N__15455),
            .I(\Inst_eia232.Inst_receiver.n5597_cascade_ ));
    InMux I__1848 (
            .O(N__15452),
            .I(N__15449));
    LocalMux I__1847 (
            .O(N__15449),
            .I(\Inst_eia232.xoff ));
    CascadeMux I__1846 (
            .O(N__15446),
            .I(\Inst_eia232.Inst_receiver.n90_cascade_ ));
    CascadeMux I__1845 (
            .O(N__15443),
            .I(\Inst_eia232.Inst_receiver.n8831_cascade_ ));
    CEMux I__1844 (
            .O(N__15440),
            .I(N__15437));
    LocalMux I__1843 (
            .O(N__15437),
            .I(N__15434));
    Span4Mux_h I__1842 (
            .O(N__15434),
            .I(N__15431));
    Odrv4 I__1841 (
            .O(N__15431),
            .I(\Inst_eia232.Inst_transmitter.n3552 ));
    CascadeMux I__1840 (
            .O(N__15428),
            .I(\Inst_eia232.Inst_receiver.n7_adj_1264_cascade_ ));
    CascadeMux I__1839 (
            .O(N__15425),
            .I(\Inst_eia232.Inst_receiver.n8769_cascade_ ));
    CascadeMux I__1838 (
            .O(N__15422),
            .I(\Inst_eia232.Inst_receiver.n6736_cascade_ ));
    InMux I__1837 (
            .O(N__15419),
            .I(N__15416));
    LocalMux I__1836 (
            .O(N__15416),
            .I(\Inst_eia232.Inst_receiver.n8772 ));
    InMux I__1835 (
            .O(N__15413),
            .I(N__15401));
    InMux I__1834 (
            .O(N__15412),
            .I(N__15401));
    InMux I__1833 (
            .O(N__15411),
            .I(N__15401));
    InMux I__1832 (
            .O(N__15410),
            .I(N__15401));
    LocalMux I__1831 (
            .O(N__15401),
            .I(\Inst_eia232.Inst_receiver.bytecount_2 ));
    CascadeMux I__1830 (
            .O(N__15398),
            .I(N__15392));
    InMux I__1829 (
            .O(N__15397),
            .I(N__15388));
    InMux I__1828 (
            .O(N__15396),
            .I(N__15379));
    InMux I__1827 (
            .O(N__15395),
            .I(N__15379));
    InMux I__1826 (
            .O(N__15392),
            .I(N__15379));
    InMux I__1825 (
            .O(N__15391),
            .I(N__15379));
    LocalMux I__1824 (
            .O(N__15388),
            .I(\Inst_eia232.Inst_receiver.bytecount_1 ));
    LocalMux I__1823 (
            .O(N__15379),
            .I(\Inst_eia232.Inst_receiver.bytecount_1 ));
    CascadeMux I__1822 (
            .O(N__15374),
            .I(\Inst_eia232.Inst_receiver.n8582_cascade_ ));
    InMux I__1821 (
            .O(N__15371),
            .I(N__15368));
    LocalMux I__1820 (
            .O(N__15368),
            .I(\GENERIC_FIFO_1.n18_adj_1277 ));
    CascadeMux I__1819 (
            .O(N__15365),
            .I(\GENERIC_FIFO_1.n141_cascade_ ));
    CascadeMux I__1818 (
            .O(N__15362),
            .I(N__15359));
    CascadeBuf I__1817 (
            .O(N__15359),
            .I(N__15356));
    CascadeMux I__1816 (
            .O(N__15356),
            .I(N__15353));
    InMux I__1815 (
            .O(N__15353),
            .I(N__15350));
    LocalMux I__1814 (
            .O(N__15350),
            .I(N__15347));
    Span4Mux_h I__1813 (
            .O(N__15347),
            .I(N__15344));
    Odrv4 I__1812 (
            .O(N__15344),
            .I(\GENERIC_FIFO_1.n69 ));
    CascadeMux I__1811 (
            .O(N__15341),
            .I(\Inst_eia232.Inst_receiver.n2143_cascade_ ));
    CascadeMux I__1810 (
            .O(N__15338),
            .I(N__15333));
    InMux I__1809 (
            .O(N__15337),
            .I(N__15323));
    InMux I__1808 (
            .O(N__15336),
            .I(N__15323));
    InMux I__1807 (
            .O(N__15333),
            .I(N__15323));
    InMux I__1806 (
            .O(N__15332),
            .I(N__15323));
    LocalMux I__1805 (
            .O(N__15323),
            .I(\Inst_eia232.Inst_receiver.bitcount_1 ));
    CascadeMux I__1804 (
            .O(N__15320),
            .I(N__15316));
    InMux I__1803 (
            .O(N__15319),
            .I(N__15308));
    InMux I__1802 (
            .O(N__15316),
            .I(N__15308));
    InMux I__1801 (
            .O(N__15315),
            .I(N__15308));
    LocalMux I__1800 (
            .O(N__15308),
            .I(\Inst_eia232.Inst_receiver.bitcount_2 ));
    CascadeMux I__1799 (
            .O(N__15305),
            .I(N__15301));
    InMux I__1798 (
            .O(N__15304),
            .I(N__15296));
    InMux I__1797 (
            .O(N__15301),
            .I(N__15296));
    LocalMux I__1796 (
            .O(N__15296),
            .I(\Inst_eia232.Inst_receiver.bitcount_3 ));
    InMux I__1795 (
            .O(N__15293),
            .I(N__15278));
    InMux I__1794 (
            .O(N__15292),
            .I(N__15278));
    InMux I__1793 (
            .O(N__15291),
            .I(N__15278));
    InMux I__1792 (
            .O(N__15290),
            .I(N__15278));
    InMux I__1791 (
            .O(N__15289),
            .I(N__15278));
    LocalMux I__1790 (
            .O(N__15278),
            .I(\Inst_eia232.Inst_receiver.bitcount_0 ));
    InMux I__1789 (
            .O(N__15275),
            .I(N__15272));
    LocalMux I__1788 (
            .O(N__15272),
            .I(\GENERIC_FIFO_1.n8650 ));
    InMux I__1787 (
            .O(N__15269),
            .I(N__15266));
    LocalMux I__1786 (
            .O(N__15266),
            .I(N__15263));
    Span4Mux_s2_h I__1785 (
            .O(N__15263),
            .I(N__15260));
    Odrv4 I__1784 (
            .O(N__15260),
            .I(\GENERIC_FIFO_1.n8681 ));
    CascadeMux I__1783 (
            .O(N__15257),
            .I(N__15254));
    CascadeBuf I__1782 (
            .O(N__15254),
            .I(N__15251));
    CascadeMux I__1781 (
            .O(N__15251),
            .I(N__15248));
    InMux I__1780 (
            .O(N__15248),
            .I(N__15245));
    LocalMux I__1779 (
            .O(N__15245),
            .I(N__15242));
    Odrv4 I__1778 (
            .O(N__15242),
            .I(\GENERIC_FIFO_1.n78 ));
    CascadeMux I__1777 (
            .O(N__15239),
            .I(N__15236));
    InMux I__1776 (
            .O(N__15236),
            .I(N__15233));
    LocalMux I__1775 (
            .O(N__15233),
            .I(\GENERIC_FIFO_1.level_9__N_900 ));
    CascadeMux I__1774 (
            .O(N__15230),
            .I(N__15227));
    InMux I__1773 (
            .O(N__15227),
            .I(N__15224));
    LocalMux I__1772 (
            .O(N__15224),
            .I(N__15221));
    Odrv4 I__1771 (
            .O(N__15221),
            .I(\GENERIC_FIFO_1.n8654 ));
    InMux I__1770 (
            .O(N__15218),
            .I(N__15215));
    LocalMux I__1769 (
            .O(N__15215),
            .I(\GENERIC_FIFO_1.n1418 ));
    InMux I__1768 (
            .O(N__15212),
            .I(N__15209));
    LocalMux I__1767 (
            .O(N__15209),
            .I(N__15206));
    Odrv4 I__1766 (
            .O(N__15206),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_6 ));
    InMux I__1765 (
            .O(N__15203),
            .I(N__15200));
    LocalMux I__1764 (
            .O(N__15200),
            .I(N__15196));
    InMux I__1763 (
            .O(N__15199),
            .I(N__15193));
    Odrv4 I__1762 (
            .O(N__15196),
            .I(\GENERIC_FIFO_1.level_9_N_876_2 ));
    LocalMux I__1761 (
            .O(N__15193),
            .I(\GENERIC_FIFO_1.level_9_N_876_2 ));
    CascadeMux I__1760 (
            .O(N__15188),
            .I(N__15184));
    InMux I__1759 (
            .O(N__15187),
            .I(N__15181));
    InMux I__1758 (
            .O(N__15184),
            .I(N__15178));
    LocalMux I__1757 (
            .O(N__15181),
            .I(N__15175));
    LocalMux I__1756 (
            .O(N__15178),
            .I(\GENERIC_FIFO_1.level_9_N_876_6 ));
    Odrv4 I__1755 (
            .O(N__15175),
            .I(\GENERIC_FIFO_1.level_9_N_876_6 ));
    CascadeMux I__1754 (
            .O(N__15170),
            .I(N__15167));
    InMux I__1753 (
            .O(N__15167),
            .I(N__15164));
    LocalMux I__1752 (
            .O(N__15164),
            .I(N__15160));
    InMux I__1751 (
            .O(N__15163),
            .I(N__15157));
    Odrv4 I__1750 (
            .O(N__15160),
            .I(\GENERIC_FIFO_1.level_9_N_876_0 ));
    LocalMux I__1749 (
            .O(N__15157),
            .I(\GENERIC_FIFO_1.level_9_N_876_0 ));
    InMux I__1748 (
            .O(N__15152),
            .I(N__15148));
    InMux I__1747 (
            .O(N__15151),
            .I(N__15145));
    LocalMux I__1746 (
            .O(N__15148),
            .I(\GENERIC_FIFO_1.level_9_N_876_8 ));
    LocalMux I__1745 (
            .O(N__15145),
            .I(\GENERIC_FIFO_1.level_9_N_876_8 ));
    InMux I__1744 (
            .O(N__15140),
            .I(N__15137));
    LocalMux I__1743 (
            .O(N__15137),
            .I(N__15133));
    InMux I__1742 (
            .O(N__15136),
            .I(N__15130));
    Odrv4 I__1741 (
            .O(N__15133),
            .I(\GENERIC_FIFO_1.level_9_N_876_5 ));
    LocalMux I__1740 (
            .O(N__15130),
            .I(\GENERIC_FIFO_1.level_9_N_876_5 ));
    CascadeMux I__1739 (
            .O(N__15125),
            .I(\GENERIC_FIFO_1.n16_adj_1276_cascade_ ));
    InMux I__1738 (
            .O(N__15122),
            .I(N__15118));
    InMux I__1737 (
            .O(N__15121),
            .I(N__15115));
    LocalMux I__1736 (
            .O(N__15118),
            .I(\GENERIC_FIFO_1.level_9_N_876_9 ));
    LocalMux I__1735 (
            .O(N__15115),
            .I(\GENERIC_FIFO_1.level_9_N_876_9 ));
    InMux I__1734 (
            .O(N__15110),
            .I(N__15107));
    LocalMux I__1733 (
            .O(N__15107),
            .I(\GENERIC_FIFO_1.n17_adj_1278 ));
    CascadeMux I__1732 (
            .O(N__15104),
            .I(N__15101));
    InMux I__1731 (
            .O(N__15101),
            .I(N__15098));
    LocalMux I__1730 (
            .O(N__15098),
            .I(N__15095));
    Odrv12 I__1729 (
            .O(N__15095),
            .I(\GENERIC_FIFO_1.n1396 ));
    CascadeMux I__1728 (
            .O(N__15092),
            .I(N__15089));
    InMux I__1727 (
            .O(N__15089),
            .I(N__15086));
    LocalMux I__1726 (
            .O(N__15086),
            .I(\GENERIC_FIFO_1.n22 ));
    InMux I__1725 (
            .O(N__15083),
            .I(\GENERIC_FIFO_1.n7810 ));
    CascadeMux I__1724 (
            .O(N__15080),
            .I(N__15077));
    InMux I__1723 (
            .O(N__15077),
            .I(N__15074));
    LocalMux I__1722 (
            .O(N__15074),
            .I(\GENERIC_FIFO_1.n21 ));
    InMux I__1721 (
            .O(N__15071),
            .I(\GENERIC_FIFO_1.n7811 ));
    CascadeMux I__1720 (
            .O(N__15068),
            .I(N__15065));
    InMux I__1719 (
            .O(N__15065),
            .I(N__15062));
    LocalMux I__1718 (
            .O(N__15062),
            .I(\GENERIC_FIFO_1.n20 ));
    InMux I__1717 (
            .O(N__15059),
            .I(\GENERIC_FIFO_1.n7812 ));
    CascadeMux I__1716 (
            .O(N__15056),
            .I(N__15053));
    InMux I__1715 (
            .O(N__15053),
            .I(N__15050));
    LocalMux I__1714 (
            .O(N__15050),
            .I(\GENERIC_FIFO_1.n19 ));
    InMux I__1713 (
            .O(N__15047),
            .I(\GENERIC_FIFO_1.n7813 ));
    CascadeMux I__1712 (
            .O(N__15044),
            .I(N__15041));
    InMux I__1711 (
            .O(N__15041),
            .I(N__15038));
    LocalMux I__1710 (
            .O(N__15038),
            .I(N__15035));
    Odrv4 I__1709 (
            .O(N__15035),
            .I(\GENERIC_FIFO_1.n18_adj_1275 ));
    InMux I__1708 (
            .O(N__15032),
            .I(\GENERIC_FIFO_1.n7814 ));
    CascadeMux I__1707 (
            .O(N__15029),
            .I(N__15026));
    InMux I__1706 (
            .O(N__15026),
            .I(N__15023));
    LocalMux I__1705 (
            .O(N__15023),
            .I(\GENERIC_FIFO_1.n17 ));
    InMux I__1704 (
            .O(N__15020),
            .I(\GENERIC_FIFO_1.n7815 ));
    InMux I__1703 (
            .O(N__15017),
            .I(N__15014));
    LocalMux I__1702 (
            .O(N__15014),
            .I(\GENERIC_FIFO_1.n16_adj_1273 ));
    InMux I__1701 (
            .O(N__15011),
            .I(bfn_2_14_0_));
    InMux I__1700 (
            .O(N__15008),
            .I(\GENERIC_FIFO_1.n7817 ));
    InMux I__1699 (
            .O(N__15005),
            .I(N__15002));
    LocalMux I__1698 (
            .O(N__15002),
            .I(\GENERIC_FIFO_1.n15 ));
    CascadeMux I__1697 (
            .O(N__14999),
            .I(\GENERIC_FIFO_1.n18_cascade_ ));
    CEMux I__1696 (
            .O(N__14996),
            .I(N__14993));
    LocalMux I__1695 (
            .O(N__14993),
            .I(N__14988));
    SRMux I__1694 (
            .O(N__14992),
            .I(N__14985));
    SRMux I__1693 (
            .O(N__14991),
            .I(N__14982));
    Span4Mux_v I__1692 (
            .O(N__14988),
            .I(N__14978));
    LocalMux I__1691 (
            .O(N__14985),
            .I(N__14975));
    LocalMux I__1690 (
            .O(N__14982),
            .I(N__14972));
    CEMux I__1689 (
            .O(N__14981),
            .I(N__14968));
    Span4Mux_s1_h I__1688 (
            .O(N__14978),
            .I(N__14963));
    Span4Mux_h I__1687 (
            .O(N__14975),
            .I(N__14963));
    Span4Mux_h I__1686 (
            .O(N__14972),
            .I(N__14960));
    InMux I__1685 (
            .O(N__14971),
            .I(N__14957));
    LocalMux I__1684 (
            .O(N__14968),
            .I(\GENERIC_FIFO_1.fifo_memory_N_983 ));
    Odrv4 I__1683 (
            .O(N__14963),
            .I(\GENERIC_FIFO_1.fifo_memory_N_983 ));
    Odrv4 I__1682 (
            .O(N__14960),
            .I(\GENERIC_FIFO_1.fifo_memory_N_983 ));
    LocalMux I__1681 (
            .O(N__14957),
            .I(\GENERIC_FIFO_1.fifo_memory_N_983 ));
    CascadeMux I__1680 (
            .O(N__14948),
            .I(N__14945));
    CascadeBuf I__1679 (
            .O(N__14945),
            .I(N__14942));
    CascadeMux I__1678 (
            .O(N__14942),
            .I(N__14939));
    InMux I__1677 (
            .O(N__14939),
            .I(N__14935));
    InMux I__1676 (
            .O(N__14938),
            .I(N__14931));
    LocalMux I__1675 (
            .O(N__14935),
            .I(N__14926));
    InMux I__1674 (
            .O(N__14934),
            .I(N__14923));
    LocalMux I__1673 (
            .O(N__14931),
            .I(N__14920));
    InMux I__1672 (
            .O(N__14930),
            .I(N__14915));
    InMux I__1671 (
            .O(N__14929),
            .I(N__14915));
    Span4Mux_h I__1670 (
            .O(N__14926),
            .I(N__14912));
    LocalMux I__1669 (
            .O(N__14923),
            .I(\GENERIC_FIFO_1.write_pointer_4 ));
    Odrv12 I__1668 (
            .O(N__14920),
            .I(\GENERIC_FIFO_1.write_pointer_4 ));
    LocalMux I__1667 (
            .O(N__14915),
            .I(\GENERIC_FIFO_1.write_pointer_4 ));
    Odrv4 I__1666 (
            .O(N__14912),
            .I(\GENERIC_FIFO_1.write_pointer_4 ));
    InMux I__1665 (
            .O(N__14903),
            .I(N__14900));
    LocalMux I__1664 (
            .O(N__14900),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_4 ));
    InMux I__1663 (
            .O(N__14897),
            .I(N__14894));
    LocalMux I__1662 (
            .O(N__14894),
            .I(N__14891));
    Odrv4 I__1661 (
            .O(N__14891),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_5 ));
    InMux I__1660 (
            .O(N__14888),
            .I(N__14885));
    LocalMux I__1659 (
            .O(N__14885),
            .I(N__14882));
    Odrv12 I__1658 (
            .O(N__14882),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n11 ));
    CascadeMux I__1657 (
            .O(N__14879),
            .I(N__14876));
    CascadeBuf I__1656 (
            .O(N__14876),
            .I(N__14872));
    InMux I__1655 (
            .O(N__14875),
            .I(N__14869));
    CascadeMux I__1654 (
            .O(N__14872),
            .I(N__14865));
    LocalMux I__1653 (
            .O(N__14869),
            .I(N__14860));
    InMux I__1652 (
            .O(N__14868),
            .I(N__14857));
    InMux I__1651 (
            .O(N__14865),
            .I(N__14854));
    InMux I__1650 (
            .O(N__14864),
            .I(N__14851));
    InMux I__1649 (
            .O(N__14863),
            .I(N__14848));
    Span4Mux_s2_v I__1648 (
            .O(N__14860),
            .I(N__14843));
    LocalMux I__1647 (
            .O(N__14857),
            .I(N__14843));
    LocalMux I__1646 (
            .O(N__14854),
            .I(N__14840));
    LocalMux I__1645 (
            .O(N__14851),
            .I(\GENERIC_FIFO_1.write_pointer_5 ));
    LocalMux I__1644 (
            .O(N__14848),
            .I(\GENERIC_FIFO_1.write_pointer_5 ));
    Odrv4 I__1643 (
            .O(N__14843),
            .I(\GENERIC_FIFO_1.write_pointer_5 ));
    Odrv12 I__1642 (
            .O(N__14840),
            .I(\GENERIC_FIFO_1.write_pointer_5 ));
    CascadeMux I__1641 (
            .O(N__14831),
            .I(\GENERIC_FIFO_1.n16_cascade_ ));
    InMux I__1640 (
            .O(N__14828),
            .I(N__14825));
    LocalMux I__1639 (
            .O(N__14825),
            .I(\GENERIC_FIFO_1.n20_adj_1274 ));
    SRMux I__1638 (
            .O(N__14822),
            .I(N__14818));
    SRMux I__1637 (
            .O(N__14821),
            .I(N__14815));
    LocalMux I__1636 (
            .O(N__14818),
            .I(\GENERIC_FIFO_1.n4721 ));
    LocalMux I__1635 (
            .O(N__14815),
            .I(\GENERIC_FIFO_1.n4721 ));
    InMux I__1634 (
            .O(N__14810),
            .I(N__14807));
    LocalMux I__1633 (
            .O(N__14807),
            .I(N__14804));
    Odrv4 I__1632 (
            .O(N__14804),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9105 ));
    InMux I__1631 (
            .O(N__14801),
            .I(N__14798));
    LocalMux I__1630 (
            .O(N__14798),
            .I(N__14795));
    Odrv12 I__1629 (
            .O(N__14795),
            .I(\GENERIC_FIFO_1.level_9_N_925_0 ));
    InMux I__1628 (
            .O(N__14792),
            .I(N__14789));
    LocalMux I__1627 (
            .O(N__14789),
            .I(\GENERIC_FIFO_1.n24 ));
    CascadeMux I__1626 (
            .O(N__14786),
            .I(N__14783));
    InMux I__1625 (
            .O(N__14783),
            .I(N__14780));
    LocalMux I__1624 (
            .O(N__14780),
            .I(\GENERIC_FIFO_1.n23 ));
    InMux I__1623 (
            .O(N__14777),
            .I(\GENERIC_FIFO_1.n7809 ));
    InMux I__1622 (
            .O(N__14774),
            .I(N__14770));
    InMux I__1621 (
            .O(N__14773),
            .I(N__14767));
    LocalMux I__1620 (
            .O(N__14770),
            .I(N__14764));
    LocalMux I__1619 (
            .O(N__14767),
            .I(maskRegister_5));
    Odrv4 I__1618 (
            .O(N__14764),
            .I(maskRegister_5));
    InMux I__1617 (
            .O(N__14759),
            .I(N__14755));
    InMux I__1616 (
            .O(N__14758),
            .I(N__14746));
    LocalMux I__1615 (
            .O(N__14755),
            .I(N__14743));
    InMux I__1614 (
            .O(N__14754),
            .I(N__14738));
    InMux I__1613 (
            .O(N__14753),
            .I(N__14738));
    InMux I__1612 (
            .O(N__14752),
            .I(N__14729));
    InMux I__1611 (
            .O(N__14751),
            .I(N__14729));
    InMux I__1610 (
            .O(N__14750),
            .I(N__14729));
    InMux I__1609 (
            .O(N__14749),
            .I(N__14729));
    LocalMux I__1608 (
            .O(N__14746),
            .I(N__14724));
    Span4Mux_v I__1607 (
            .O(N__14743),
            .I(N__14724));
    LocalMux I__1606 (
            .O(N__14738),
            .I(\Inst_eia232.Inst_transmitter.n6703 ));
    LocalMux I__1605 (
            .O(N__14729),
            .I(\Inst_eia232.Inst_transmitter.n6703 ));
    Odrv4 I__1604 (
            .O(N__14724),
            .I(\Inst_eia232.Inst_transmitter.n6703 ));
    CascadeMux I__1603 (
            .O(N__14717),
            .I(N__14714));
    InMux I__1602 (
            .O(N__14714),
            .I(N__14711));
    LocalMux I__1601 (
            .O(N__14711),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_5 ));
    InMux I__1600 (
            .O(N__14708),
            .I(N__14705));
    LocalMux I__1599 (
            .O(N__14705),
            .I(N__14702));
    Span4Mux_v I__1598 (
            .O(N__14702),
            .I(N__14698));
    InMux I__1597 (
            .O(N__14701),
            .I(N__14695));
    Odrv4 I__1596 (
            .O(N__14698),
            .I(\Inst_eia232.Inst_transmitter.byte_5 ));
    LocalMux I__1595 (
            .O(N__14695),
            .I(\Inst_eia232.Inst_transmitter.byte_5 ));
    CascadeMux I__1594 (
            .O(N__14690),
            .I(\GENERIC_FIFO_1.n8677_cascade_ ));
    CascadeMux I__1593 (
            .O(N__14687),
            .I(\GENERIC_FIFO_1.n1396_cascade_ ));
    SRMux I__1592 (
            .O(N__14684),
            .I(N__14681));
    LocalMux I__1591 (
            .O(N__14681),
            .I(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4743 ));
    InMux I__1590 (
            .O(N__14678),
            .I(N__14675));
    LocalMux I__1589 (
            .O(N__14675),
            .I(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_0 ));
    CascadeMux I__1588 (
            .O(N__14672),
            .I(N__14669));
    CascadeBuf I__1587 (
            .O(N__14669),
            .I(N__14666));
    CascadeMux I__1586 (
            .O(N__14666),
            .I(N__14663));
    InMux I__1585 (
            .O(N__14663),
            .I(N__14658));
    InMux I__1584 (
            .O(N__14662),
            .I(N__14651));
    InMux I__1583 (
            .O(N__14661),
            .I(N__14651));
    LocalMux I__1582 (
            .O(N__14658),
            .I(N__14648));
    InMux I__1581 (
            .O(N__14657),
            .I(N__14645));
    InMux I__1580 (
            .O(N__14656),
            .I(N__14642));
    LocalMux I__1579 (
            .O(N__14651),
            .I(N__14639));
    Span4Mux_v I__1578 (
            .O(N__14648),
            .I(N__14636));
    LocalMux I__1577 (
            .O(N__14645),
            .I(\GENERIC_FIFO_1.write_pointer_8 ));
    LocalMux I__1576 (
            .O(N__14642),
            .I(\GENERIC_FIFO_1.write_pointer_8 ));
    Odrv12 I__1575 (
            .O(N__14639),
            .I(\GENERIC_FIFO_1.write_pointer_8 ));
    Odrv4 I__1574 (
            .O(N__14636),
            .I(\GENERIC_FIFO_1.write_pointer_8 ));
    CascadeMux I__1573 (
            .O(N__14627),
            .I(N__14624));
    CascadeBuf I__1572 (
            .O(N__14624),
            .I(N__14621));
    CascadeMux I__1571 (
            .O(N__14621),
            .I(N__14618));
    InMux I__1570 (
            .O(N__14618),
            .I(N__14612));
    CascadeMux I__1569 (
            .O(N__14617),
            .I(N__14608));
    InMux I__1568 (
            .O(N__14616),
            .I(N__14603));
    InMux I__1567 (
            .O(N__14615),
            .I(N__14603));
    LocalMux I__1566 (
            .O(N__14612),
            .I(N__14600));
    InMux I__1565 (
            .O(N__14611),
            .I(N__14597));
    InMux I__1564 (
            .O(N__14608),
            .I(N__14594));
    LocalMux I__1563 (
            .O(N__14603),
            .I(N__14591));
    Span4Mux_v I__1562 (
            .O(N__14600),
            .I(N__14588));
    LocalMux I__1561 (
            .O(N__14597),
            .I(\GENERIC_FIFO_1.write_pointer_9 ));
    LocalMux I__1560 (
            .O(N__14594),
            .I(\GENERIC_FIFO_1.write_pointer_9 ));
    Odrv12 I__1559 (
            .O(N__14591),
            .I(\GENERIC_FIFO_1.write_pointer_9 ));
    Odrv4 I__1558 (
            .O(N__14588),
            .I(\GENERIC_FIFO_1.write_pointer_9 ));
    CascadeMux I__1557 (
            .O(N__14579),
            .I(N__14576));
    CascadeBuf I__1556 (
            .O(N__14576),
            .I(N__14573));
    CascadeMux I__1555 (
            .O(N__14573),
            .I(N__14568));
    InMux I__1554 (
            .O(N__14572),
            .I(N__14563));
    InMux I__1553 (
            .O(N__14571),
            .I(N__14560));
    InMux I__1552 (
            .O(N__14568),
            .I(N__14557));
    InMux I__1551 (
            .O(N__14567),
            .I(N__14554));
    InMux I__1550 (
            .O(N__14566),
            .I(N__14551));
    LocalMux I__1549 (
            .O(N__14563),
            .I(N__14546));
    LocalMux I__1548 (
            .O(N__14560),
            .I(N__14546));
    LocalMux I__1547 (
            .O(N__14557),
            .I(N__14543));
    LocalMux I__1546 (
            .O(N__14554),
            .I(\GENERIC_FIFO_1.write_pointer_7 ));
    LocalMux I__1545 (
            .O(N__14551),
            .I(\GENERIC_FIFO_1.write_pointer_7 ));
    Odrv12 I__1544 (
            .O(N__14546),
            .I(\GENERIC_FIFO_1.write_pointer_7 ));
    Odrv12 I__1543 (
            .O(N__14543),
            .I(\GENERIC_FIFO_1.write_pointer_7 ));
    InMux I__1542 (
            .O(N__14534),
            .I(\GENERIC_FIFO_1.n7930 ));
    InMux I__1541 (
            .O(N__14531),
            .I(\GENERIC_FIFO_1.n7931 ));
    InMux I__1540 (
            .O(N__14528),
            .I(\GENERIC_FIFO_1.n7932 ));
    InMux I__1539 (
            .O(N__14525),
            .I(\GENERIC_FIFO_1.n7933 ));
    InMux I__1538 (
            .O(N__14522),
            .I(\GENERIC_FIFO_1.n7934 ));
    InMux I__1537 (
            .O(N__14519),
            .I(\GENERIC_FIFO_1.n7935 ));
    InMux I__1536 (
            .O(N__14516),
            .I(bfn_2_9_0_));
    InMux I__1535 (
            .O(N__14513),
            .I(\GENERIC_FIFO_1.n7937 ));
    InMux I__1534 (
            .O(N__14510),
            .I(N__14504));
    InMux I__1533 (
            .O(N__14509),
            .I(N__14504));
    LocalMux I__1532 (
            .O(N__14504),
            .I(disabledGroupsReg_3));
    InMux I__1531 (
            .O(N__14501),
            .I(N__14497));
    InMux I__1530 (
            .O(N__14500),
            .I(N__14494));
    LocalMux I__1529 (
            .O(N__14497),
            .I(N__14491));
    LocalMux I__1528 (
            .O(N__14494),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_2 ));
    Odrv4 I__1527 (
            .O(N__14491),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_2 ));
    CascadeMux I__1526 (
            .O(N__14486),
            .I(N__14483));
    InMux I__1525 (
            .O(N__14483),
            .I(N__14477));
    InMux I__1524 (
            .O(N__14482),
            .I(N__14477));
    LocalMux I__1523 (
            .O(N__14477),
            .I(disabledGroupsReg_2));
    InMux I__1522 (
            .O(N__14474),
            .I(N__14471));
    LocalMux I__1521 (
            .O(N__14471),
            .I(N__14468));
    Span4Mux_s2_h I__1520 (
            .O(N__14468),
            .I(N__14464));
    InMux I__1519 (
            .O(N__14467),
            .I(N__14461));
    Odrv4 I__1518 (
            .O(N__14464),
            .I(\Inst_eia232.Inst_transmitter.byte_7 ));
    LocalMux I__1517 (
            .O(N__14461),
            .I(\Inst_eia232.Inst_transmitter.byte_7 ));
    InMux I__1516 (
            .O(N__14456),
            .I(N__14453));
    LocalMux I__1515 (
            .O(N__14453),
            .I(N__14450));
    Span4Mux_v I__1514 (
            .O(N__14450),
            .I(N__14447));
    Odrv4 I__1513 (
            .O(N__14447),
            .I(outputdata_7));
    CascadeMux I__1512 (
            .O(N__14444),
            .I(N__14440));
    CascadeMux I__1511 (
            .O(N__14443),
            .I(N__14437));
    InMux I__1510 (
            .O(N__14440),
            .I(N__14432));
    InMux I__1509 (
            .O(N__14437),
            .I(N__14432));
    LocalMux I__1508 (
            .O(N__14432),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_7 ));
    InMux I__1507 (
            .O(N__14429),
            .I(bfn_2_8_0_));
    InMux I__1506 (
            .O(N__14426),
            .I(\GENERIC_FIFO_1.n7929 ));
    CascadeMux I__1505 (
            .O(N__14423),
            .I(N__14419));
    InMux I__1504 (
            .O(N__14422),
            .I(N__14405));
    InMux I__1503 (
            .O(N__14419),
            .I(N__14405));
    InMux I__1502 (
            .O(N__14418),
            .I(N__14405));
    InMux I__1501 (
            .O(N__14417),
            .I(N__14400));
    InMux I__1500 (
            .O(N__14416),
            .I(N__14400));
    InMux I__1499 (
            .O(N__14415),
            .I(N__14391));
    InMux I__1498 (
            .O(N__14414),
            .I(N__14391));
    InMux I__1497 (
            .O(N__14413),
            .I(N__14391));
    InMux I__1496 (
            .O(N__14412),
            .I(N__14391));
    LocalMux I__1495 (
            .O(N__14405),
            .I(bytes_0));
    LocalMux I__1494 (
            .O(N__14400),
            .I(bytes_0));
    LocalMux I__1493 (
            .O(N__14391),
            .I(bytes_0));
    CascadeMux I__1492 (
            .O(N__14384),
            .I(\Inst_eia232.Inst_transmitter.n3652_cascade_ ));
    InMux I__1491 (
            .O(N__14381),
            .I(N__14378));
    LocalMux I__1490 (
            .O(N__14378),
            .I(n1336));
    InMux I__1489 (
            .O(N__14375),
            .I(N__14372));
    LocalMux I__1488 (
            .O(N__14372),
            .I(N__14369));
    Span4Mux_v I__1487 (
            .O(N__14369),
            .I(N__14366));
    Odrv4 I__1486 (
            .O(N__14366),
            .I(outputdata_1));
    CascadeMux I__1485 (
            .O(N__14363),
            .I(N__14359));
    InMux I__1484 (
            .O(N__14362),
            .I(N__14356));
    InMux I__1483 (
            .O(N__14359),
            .I(N__14353));
    LocalMux I__1482 (
            .O(N__14356),
            .I(N__14350));
    LocalMux I__1481 (
            .O(N__14353),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_1 ));
    Odrv12 I__1480 (
            .O(N__14350),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_1 ));
    InMux I__1479 (
            .O(N__14345),
            .I(N__14342));
    LocalMux I__1478 (
            .O(N__14342),
            .I(N__14339));
    Sp12to4 I__1477 (
            .O(N__14339),
            .I(N__14336));
    Odrv12 I__1476 (
            .O(N__14336),
            .I(outputdata_2));
    InMux I__1475 (
            .O(N__14333),
            .I(N__14329));
    InMux I__1474 (
            .O(N__14332),
            .I(N__14326));
    LocalMux I__1473 (
            .O(N__14329),
            .I(N__14323));
    LocalMux I__1472 (
            .O(N__14326),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_2 ));
    Odrv4 I__1471 (
            .O(N__14323),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_2 ));
    CascadeMux I__1470 (
            .O(N__14318),
            .I(N__14315));
    InMux I__1469 (
            .O(N__14315),
            .I(N__14312));
    LocalMux I__1468 (
            .O(N__14312),
            .I(N__14309));
    Span12Mux_s11_v I__1467 (
            .O(N__14309),
            .I(N__14306));
    Odrv12 I__1466 (
            .O(N__14306),
            .I(outputdata_3));
    InMux I__1465 (
            .O(N__14303),
            .I(N__14299));
    InMux I__1464 (
            .O(N__14302),
            .I(N__14296));
    LocalMux I__1463 (
            .O(N__14299),
            .I(N__14293));
    LocalMux I__1462 (
            .O(N__14296),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_3 ));
    Odrv4 I__1461 (
            .O(N__14293),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_3 ));
    InMux I__1460 (
            .O(N__14288),
            .I(N__14285));
    LocalMux I__1459 (
            .O(N__14285),
            .I(N__14282));
    Span4Mux_s2_h I__1458 (
            .O(N__14282),
            .I(N__14279));
    Odrv4 I__1457 (
            .O(N__14279),
            .I(outputdata_6));
    InMux I__1456 (
            .O(N__14276),
            .I(N__14272));
    InMux I__1455 (
            .O(N__14275),
            .I(N__14269));
    LocalMux I__1454 (
            .O(N__14272),
            .I(N__14266));
    LocalMux I__1453 (
            .O(N__14269),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_6 ));
    Odrv4 I__1452 (
            .O(N__14266),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_6 ));
    InMux I__1451 (
            .O(N__14261),
            .I(N__14257));
    InMux I__1450 (
            .O(N__14260),
            .I(N__14254));
    LocalMux I__1449 (
            .O(N__14257),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_1 ));
    LocalMux I__1448 (
            .O(N__14254),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_1 ));
    InMux I__1447 (
            .O(N__14249),
            .I(N__14243));
    InMux I__1446 (
            .O(N__14248),
            .I(N__14243));
    LocalMux I__1445 (
            .O(N__14243),
            .I(disabledGroupsReg_1));
    InMux I__1444 (
            .O(N__14240),
            .I(N__14236));
    InMux I__1443 (
            .O(N__14239),
            .I(N__14233));
    LocalMux I__1442 (
            .O(N__14236),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_3 ));
    LocalMux I__1441 (
            .O(N__14233),
            .I(\Inst_eia232.Inst_transmitter.disabledBuffer_3 ));
    CascadeMux I__1440 (
            .O(N__14228),
            .I(n1320_cascade_));
    InMux I__1439 (
            .O(N__14225),
            .I(N__14221));
    InMux I__1438 (
            .O(N__14224),
            .I(N__14218));
    LocalMux I__1437 (
            .O(N__14221),
            .I(dataBuffer_28));
    LocalMux I__1436 (
            .O(N__14218),
            .I(dataBuffer_28));
    CascadeMux I__1435 (
            .O(N__14213),
            .I(\Inst_eia232.Inst_transmitter.n8756_cascade_ ));
    InMux I__1434 (
            .O(N__14210),
            .I(N__14207));
    LocalMux I__1433 (
            .O(N__14207),
            .I(N__14204));
    Span4Mux_v I__1432 (
            .O(N__14204),
            .I(N__14201));
    Span4Mux_h I__1431 (
            .O(N__14201),
            .I(N__14198));
    Odrv4 I__1430 (
            .O(N__14198),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_4 ));
    InMux I__1429 (
            .O(N__14195),
            .I(N__14192));
    LocalMux I__1428 (
            .O(N__14192),
            .I(\Inst_eia232.Inst_transmitter.byte_4 ));
    CascadeMux I__1427 (
            .O(N__14189),
            .I(state_1_N_371_1_cascade_));
    InMux I__1426 (
            .O(N__14186),
            .I(N__14183));
    LocalMux I__1425 (
            .O(N__14183),
            .I(\Inst_eia232.Inst_transmitter.n1 ));
    InMux I__1424 (
            .O(N__14180),
            .I(N__14166));
    InMux I__1423 (
            .O(N__14179),
            .I(N__14166));
    InMux I__1422 (
            .O(N__14178),
            .I(N__14166));
    InMux I__1421 (
            .O(N__14177),
            .I(N__14161));
    InMux I__1420 (
            .O(N__14176),
            .I(N__14161));
    InMux I__1419 (
            .O(N__14175),
            .I(N__14154));
    InMux I__1418 (
            .O(N__14174),
            .I(N__14154));
    InMux I__1417 (
            .O(N__14173),
            .I(N__14154));
    LocalMux I__1416 (
            .O(N__14166),
            .I(bytes_1));
    LocalMux I__1415 (
            .O(N__14161),
            .I(bytes_1));
    LocalMux I__1414 (
            .O(N__14154),
            .I(bytes_1));
    InMux I__1413 (
            .O(N__14147),
            .I(N__14137));
    InMux I__1412 (
            .O(N__14146),
            .I(N__14137));
    InMux I__1411 (
            .O(N__14145),
            .I(N__14134));
    InMux I__1410 (
            .O(N__14144),
            .I(N__14131));
    InMux I__1409 (
            .O(N__14143),
            .I(N__14126));
    InMux I__1408 (
            .O(N__14142),
            .I(N__14126));
    LocalMux I__1407 (
            .O(N__14137),
            .I(bytes_2));
    LocalMux I__1406 (
            .O(N__14134),
            .I(bytes_2));
    LocalMux I__1405 (
            .O(N__14131),
            .I(bytes_2));
    LocalMux I__1404 (
            .O(N__14126),
            .I(bytes_2));
    CascadeMux I__1403 (
            .O(N__14117),
            .I(\Inst_eia232.Inst_transmitter.n9218_cascade_ ));
    InMux I__1402 (
            .O(N__14114),
            .I(N__14111));
    LocalMux I__1401 (
            .O(N__14111),
            .I(\Inst_eia232.Inst_transmitter.n3 ));
    InMux I__1400 (
            .O(N__14108),
            .I(N__14105));
    LocalMux I__1399 (
            .O(N__14105),
            .I(N__14102));
    Odrv4 I__1398 (
            .O(N__14102),
            .I(disabled));
    CEMux I__1397 (
            .O(N__14099),
            .I(N__14096));
    LocalMux I__1396 (
            .O(N__14096),
            .I(N__14093));
    Odrv4 I__1395 (
            .O(N__14093),
            .I(\Inst_eia232.Inst_transmitter.n6745 ));
    InMux I__1394 (
            .O(N__14090),
            .I(N__14083));
    InMux I__1393 (
            .O(N__14089),
            .I(N__14083));
    InMux I__1392 (
            .O(N__14088),
            .I(N__14080));
    LocalMux I__1391 (
            .O(N__14083),
            .I(state_1_N_371_1));
    LocalMux I__1390 (
            .O(N__14080),
            .I(state_1_N_371_1));
    CEMux I__1389 (
            .O(N__14075),
            .I(N__14072));
    LocalMux I__1388 (
            .O(N__14072),
            .I(N__14068));
    CEMux I__1387 (
            .O(N__14071),
            .I(N__14065));
    Span4Mux_s3_v I__1386 (
            .O(N__14068),
            .I(N__14060));
    LocalMux I__1385 (
            .O(N__14065),
            .I(N__14060));
    Span4Mux_h I__1384 (
            .O(N__14060),
            .I(N__14056));
    InMux I__1383 (
            .O(N__14059),
            .I(N__14053));
    Odrv4 I__1382 (
            .O(N__14056),
            .I(\Inst_eia232.Inst_transmitter.n3652 ));
    LocalMux I__1381 (
            .O(N__14053),
            .I(\Inst_eia232.Inst_transmitter.n3652 ));
    InMux I__1380 (
            .O(N__14048),
            .I(N__14045));
    LocalMux I__1379 (
            .O(N__14045),
            .I(\Inst_eia232.Inst_transmitter.n1323 ));
    CascadeMux I__1378 (
            .O(N__14042),
            .I(\Inst_eia232.Inst_transmitter.n3632_cascade_ ));
    InMux I__1377 (
            .O(N__14039),
            .I(N__14036));
    LocalMux I__1376 (
            .O(N__14036),
            .I(\Inst_eia232.Inst_transmitter.byte_6 ));
    CascadeMux I__1375 (
            .O(N__14033),
            .I(N__14029));
    InMux I__1374 (
            .O(N__14032),
            .I(N__14026));
    InMux I__1373 (
            .O(N__14029),
            .I(N__14023));
    LocalMux I__1372 (
            .O(N__14026),
            .I(dataBuffer_18));
    LocalMux I__1371 (
            .O(N__14023),
            .I(dataBuffer_18));
    CascadeMux I__1370 (
            .O(N__14018),
            .I(\Inst_eia232.Inst_transmitter.n8851_cascade_ ));
    InMux I__1369 (
            .O(N__14015),
            .I(N__14012));
    LocalMux I__1368 (
            .O(N__14012),
            .I(N__14009));
    Odrv12 I__1367 (
            .O(N__14009),
            .I(\Inst_eia232.Inst_transmitter.byte_2 ));
    InMux I__1366 (
            .O(N__14006),
            .I(N__14003));
    LocalMux I__1365 (
            .O(N__14003),
            .I(\Inst_eia232.Inst_transmitter.byte_1 ));
    CascadeMux I__1364 (
            .O(N__14000),
            .I(n4248_cascade_));
    CascadeMux I__1363 (
            .O(N__13997),
            .I(n1336_cascade_));
    CascadeMux I__1362 (
            .O(N__13994),
            .I(N__13991));
    InMux I__1361 (
            .O(N__13991),
            .I(N__13987));
    InMux I__1360 (
            .O(N__13990),
            .I(N__13984));
    LocalMux I__1359 (
            .O(N__13987),
            .I(dataBuffer_25));
    LocalMux I__1358 (
            .O(N__13984),
            .I(dataBuffer_25));
    InMux I__1357 (
            .O(N__13979),
            .I(N__13976));
    LocalMux I__1356 (
            .O(N__13976),
            .I(\Inst_eia232.Inst_transmitter.n8847 ));
    CascadeMux I__1355 (
            .O(N__13973),
            .I(N__13970));
    InMux I__1354 (
            .O(N__13970),
            .I(N__13967));
    LocalMux I__1353 (
            .O(N__13967),
            .I(n4248));
    CascadeMux I__1352 (
            .O(N__13964),
            .I(N__13961));
    InMux I__1351 (
            .O(N__13961),
            .I(N__13954));
    InMux I__1350 (
            .O(N__13960),
            .I(N__13951));
    InMux I__1349 (
            .O(N__13959),
            .I(N__13946));
    InMux I__1348 (
            .O(N__13958),
            .I(N__13946));
    InMux I__1347 (
            .O(N__13957),
            .I(N__13943));
    LocalMux I__1346 (
            .O(N__13954),
            .I(N__13938));
    LocalMux I__1345 (
            .O(N__13951),
            .I(N__13938));
    LocalMux I__1344 (
            .O(N__13946),
            .I(n1320));
    LocalMux I__1343 (
            .O(N__13943),
            .I(n1320));
    Odrv4 I__1342 (
            .O(N__13938),
            .I(n1320));
    InMux I__1341 (
            .O(N__13931),
            .I(N__13925));
    InMux I__1340 (
            .O(N__13930),
            .I(N__13925));
    LocalMux I__1339 (
            .O(N__13925),
            .I(dataBuffer_22));
    InMux I__1338 (
            .O(N__13922),
            .I(N__13916));
    InMux I__1337 (
            .O(N__13921),
            .I(N__13916));
    LocalMux I__1336 (
            .O(N__13916),
            .I(dataBuffer_30));
    CascadeMux I__1335 (
            .O(N__13913),
            .I(N__13909));
    InMux I__1334 (
            .O(N__13912),
            .I(N__13906));
    InMux I__1333 (
            .O(N__13909),
            .I(N__13903));
    LocalMux I__1332 (
            .O(N__13906),
            .I(dataBuffer_24));
    LocalMux I__1331 (
            .O(N__13903),
            .I(dataBuffer_24));
    InMux I__1330 (
            .O(N__13898),
            .I(N__13895));
    LocalMux I__1329 (
            .O(N__13895),
            .I(N__13892));
    Odrv12 I__1328 (
            .O(N__13892),
            .I(\Inst_eia232.Inst_transmitter.byte_0 ));
    InMux I__1327 (
            .O(N__13889),
            .I(N__13886));
    LocalMux I__1326 (
            .O(N__13886),
            .I(N__13883));
    Odrv4 I__1325 (
            .O(N__13883),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_8 ));
    InMux I__1324 (
            .O(N__13880),
            .I(N__13877));
    LocalMux I__1323 (
            .O(N__13877),
            .I(N__13874));
    Span4Mux_v I__1322 (
            .O(N__13874),
            .I(N__13871));
    Odrv4 I__1321 (
            .O(N__13871),
            .I(\Inst_eia232.Inst_transmitter.dataBuffer_0 ));
    InMux I__1320 (
            .O(N__13868),
            .I(N__13865));
    LocalMux I__1319 (
            .O(N__13865),
            .I(\Inst_eia232.Inst_transmitter.n3571 ));
    InMux I__1318 (
            .O(N__13862),
            .I(N__13858));
    InMux I__1317 (
            .O(N__13861),
            .I(N__13855));
    LocalMux I__1316 (
            .O(N__13858),
            .I(dataBuffer_19));
    LocalMux I__1315 (
            .O(N__13855),
            .I(dataBuffer_19));
    CascadeMux I__1314 (
            .O(N__13850),
            .I(\Inst_eia232.Inst_transmitter.n8854_cascade_ ));
    InMux I__1313 (
            .O(N__13847),
            .I(N__13844));
    LocalMux I__1312 (
            .O(N__13844),
            .I(\Inst_eia232.Inst_transmitter.byte_3 ));
    InMux I__1311 (
            .O(N__13841),
            .I(N__13837));
    InMux I__1310 (
            .O(N__13840),
            .I(N__13834));
    LocalMux I__1309 (
            .O(N__13837),
            .I(dataBuffer_14));
    LocalMux I__1308 (
            .O(N__13834),
            .I(dataBuffer_14));
    InMux I__1307 (
            .O(N__13829),
            .I(\GENERIC_FIFO_1.n7826 ));
    InMux I__1306 (
            .O(N__13826),
            .I(N__13823));
    LocalMux I__1305 (
            .O(N__13823),
            .I(N__13820));
    Odrv4 I__1304 (
            .O(N__13820),
            .I(\GENERIC_FIFO_1.n3 ));
    CascadeMux I__1303 (
            .O(N__13817),
            .I(n4005_cascade_));
    CascadeMux I__1302 (
            .O(N__13814),
            .I(N__13811));
    InMux I__1301 (
            .O(N__13811),
            .I(N__13808));
    LocalMux I__1300 (
            .O(N__13808),
            .I(N__13805));
    Odrv4 I__1299 (
            .O(N__13805),
            .I(\GENERIC_FIFO_1.n12 ));
    InMux I__1298 (
            .O(N__13802),
            .I(N__13799));
    LocalMux I__1297 (
            .O(N__13799),
            .I(N__13796));
    Odrv4 I__1296 (
            .O(N__13796),
            .I(\GENERIC_FIFO_1.n11 ));
    InMux I__1295 (
            .O(N__13793),
            .I(\GENERIC_FIFO_1.n7818 ));
    InMux I__1294 (
            .O(N__13790),
            .I(N__13787));
    LocalMux I__1293 (
            .O(N__13787),
            .I(N__13784));
    Odrv4 I__1292 (
            .O(N__13784),
            .I(\GENERIC_FIFO_1.n10 ));
    InMux I__1291 (
            .O(N__13781),
            .I(\GENERIC_FIFO_1.n7819 ));
    InMux I__1290 (
            .O(N__13778),
            .I(N__13775));
    LocalMux I__1289 (
            .O(N__13775),
            .I(N__13772));
    Odrv4 I__1288 (
            .O(N__13772),
            .I(\GENERIC_FIFO_1.n9 ));
    InMux I__1287 (
            .O(N__13769),
            .I(\GENERIC_FIFO_1.n7820 ));
    InMux I__1286 (
            .O(N__13766),
            .I(N__13763));
    LocalMux I__1285 (
            .O(N__13763),
            .I(N__13760));
    Span4Mux_s1_h I__1284 (
            .O(N__13760),
            .I(N__13757));
    Odrv4 I__1283 (
            .O(N__13757),
            .I(\GENERIC_FIFO_1.n8 ));
    InMux I__1282 (
            .O(N__13754),
            .I(\GENERIC_FIFO_1.n7821 ));
    InMux I__1281 (
            .O(N__13751),
            .I(N__13748));
    LocalMux I__1280 (
            .O(N__13748),
            .I(N__13745));
    Odrv4 I__1279 (
            .O(N__13745),
            .I(\GENERIC_FIFO_1.n7 ));
    InMux I__1278 (
            .O(N__13742),
            .I(\GENERIC_FIFO_1.n7822 ));
    InMux I__1277 (
            .O(N__13739),
            .I(N__13736));
    LocalMux I__1276 (
            .O(N__13736),
            .I(N__13733));
    Odrv4 I__1275 (
            .O(N__13733),
            .I(\GENERIC_FIFO_1.n6 ));
    InMux I__1274 (
            .O(N__13730),
            .I(\GENERIC_FIFO_1.n7823 ));
    InMux I__1273 (
            .O(N__13727),
            .I(N__13724));
    LocalMux I__1272 (
            .O(N__13724),
            .I(N__13721));
    Odrv4 I__1271 (
            .O(N__13721),
            .I(\GENERIC_FIFO_1.n5 ));
    InMux I__1270 (
            .O(N__13718),
            .I(\GENERIC_FIFO_1.n7824 ));
    CascadeMux I__1269 (
            .O(N__13715),
            .I(N__13712));
    InMux I__1268 (
            .O(N__13712),
            .I(N__13709));
    LocalMux I__1267 (
            .O(N__13709),
            .I(N__13706));
    Odrv4 I__1266 (
            .O(N__13706),
            .I(\GENERIC_FIFO_1.n4 ));
    InMux I__1265 (
            .O(N__13703),
            .I(bfn_1_16_0_));
    InMux I__1264 (
            .O(N__13700),
            .I(\GENERIC_FIFO_1.n7830 ));
    InMux I__1263 (
            .O(N__13697),
            .I(\GENERIC_FIFO_1.n7831 ));
    InMux I__1262 (
            .O(N__13694),
            .I(\GENERIC_FIFO_1.n7832 ));
    InMux I__1261 (
            .O(N__13691),
            .I(\GENERIC_FIFO_1.n7833 ));
    InMux I__1260 (
            .O(N__13688),
            .I(bfn_1_14_0_));
    InMux I__1259 (
            .O(N__13685),
            .I(\GENERIC_FIFO_1.n7835 ));
    InMux I__1258 (
            .O(N__13682),
            .I(N__13678));
    InMux I__1257 (
            .O(N__13681),
            .I(N__13675));
    LocalMux I__1256 (
            .O(N__13678),
            .I(N__13672));
    LocalMux I__1255 (
            .O(N__13675),
            .I(\GENERIC_FIFO_1.level_9_N_876_7 ));
    Odrv4 I__1254 (
            .O(N__13672),
            .I(\GENERIC_FIFO_1.level_9_N_876_7 ));
    InMux I__1253 (
            .O(N__13667),
            .I(N__13663));
    InMux I__1252 (
            .O(N__13666),
            .I(N__13660));
    LocalMux I__1251 (
            .O(N__13663),
            .I(\GENERIC_FIFO_1.level_9_N_876_1 ));
    LocalMux I__1250 (
            .O(N__13660),
            .I(\GENERIC_FIFO_1.level_9_N_876_1 ));
    CascadeMux I__1249 (
            .O(N__13655),
            .I(N__13651));
    CascadeMux I__1248 (
            .O(N__13654),
            .I(N__13648));
    InMux I__1247 (
            .O(N__13651),
            .I(N__13645));
    InMux I__1246 (
            .O(N__13648),
            .I(N__13642));
    LocalMux I__1245 (
            .O(N__13645),
            .I(\GENERIC_FIFO_1.level_9_N_876_4 ));
    LocalMux I__1244 (
            .O(N__13642),
            .I(\GENERIC_FIFO_1.level_9_N_876_4 ));
    InMux I__1243 (
            .O(N__13637),
            .I(N__13633));
    InMux I__1242 (
            .O(N__13636),
            .I(N__13630));
    LocalMux I__1241 (
            .O(N__13633),
            .I(\GENERIC_FIFO_1.level_9_N_876_3 ));
    LocalMux I__1240 (
            .O(N__13630),
            .I(\GENERIC_FIFO_1.level_9_N_876_3 ));
    InMux I__1239 (
            .O(N__13625),
            .I(\GENERIC_FIFO_1.n7840 ));
    InMux I__1238 (
            .O(N__13622),
            .I(\GENERIC_FIFO_1.n7841 ));
    InMux I__1237 (
            .O(N__13619),
            .I(\GENERIC_FIFO_1.n7842 ));
    InMux I__1236 (
            .O(N__13616),
            .I(bfn_1_12_0_));
    InMux I__1235 (
            .O(N__13613),
            .I(\GENERIC_FIFO_1.n7844 ));
    InMux I__1234 (
            .O(N__13610),
            .I(\GENERIC_FIFO_1.n7827 ));
    InMux I__1233 (
            .O(N__13607),
            .I(\GENERIC_FIFO_1.n7828 ));
    InMux I__1232 (
            .O(N__13604),
            .I(\GENERIC_FIFO_1.n7829 ));
    InMux I__1231 (
            .O(N__13601),
            .I(N__13598));
    LocalMux I__1230 (
            .O(N__13598),
            .I(N__13595));
    Span4Mux_s3_h I__1229 (
            .O(N__13595),
            .I(N__13592));
    Odrv4 I__1228 (
            .O(N__13592),
            .I(outputdata_0));
    InMux I__1227 (
            .O(N__13589),
            .I(N__13586));
    LocalMux I__1226 (
            .O(N__13586),
            .I(N__13583));
    Odrv12 I__1225 (
            .O(N__13583),
            .I(outputdata_4));
    InMux I__1224 (
            .O(N__13580),
            .I(N__13577));
    LocalMux I__1223 (
            .O(N__13577),
            .I(N__13574));
    Odrv4 I__1222 (
            .O(N__13574),
            .I(outputdata_5));
    InMux I__1221 (
            .O(N__13571),
            .I(N__13568));
    LocalMux I__1220 (
            .O(N__13568),
            .I(N__13565));
    Span4Mux_v I__1219 (
            .O(N__13565),
            .I(N__13562));
    Odrv4 I__1218 (
            .O(N__13562),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_1 ));
    IoInMux I__1217 (
            .O(N__13559),
            .I(N__13556));
    LocalMux I__1216 (
            .O(N__13556),
            .I(N__13553));
    Span4Mux_s0_h I__1215 (
            .O(N__13553),
            .I(N__13550));
    Odrv4 I__1214 (
            .O(N__13550),
            .I(tx_c));
    InMux I__1213 (
            .O(N__13547),
            .I(bfn_1_11_0_));
    InMux I__1212 (
            .O(N__13544),
            .I(\GENERIC_FIFO_1.n7836 ));
    InMux I__1211 (
            .O(N__13541),
            .I(\GENERIC_FIFO_1.n7837 ));
    InMux I__1210 (
            .O(N__13538),
            .I(\GENERIC_FIFO_1.n7838 ));
    InMux I__1209 (
            .O(N__13535),
            .I(\GENERIC_FIFO_1.n7839 ));
    InMux I__1208 (
            .O(N__13532),
            .I(N__13525));
    InMux I__1207 (
            .O(N__13531),
            .I(N__13525));
    InMux I__1206 (
            .O(N__13530),
            .I(N__13522));
    LocalMux I__1205 (
            .O(N__13525),
            .I(\Inst_eia232.Inst_transmitter.counter_3 ));
    LocalMux I__1204 (
            .O(N__13522),
            .I(\Inst_eia232.Inst_transmitter.counter_3 ));
    CascadeMux I__1203 (
            .O(N__13517),
            .I(\Inst_eia232.Inst_transmitter.n2201_cascade_ ));
    InMux I__1202 (
            .O(N__13514),
            .I(N__13508));
    InMux I__1201 (
            .O(N__13513),
            .I(N__13508));
    LocalMux I__1200 (
            .O(N__13508),
            .I(\Inst_eia232.Inst_transmitter.counter_4 ));
    InMux I__1199 (
            .O(N__13505),
            .I(N__13502));
    LocalMux I__1198 (
            .O(N__13502),
            .I(\Inst_eia232.Inst_transmitter.n8642 ));
    InMux I__1197 (
            .O(N__13499),
            .I(N__13484));
    InMux I__1196 (
            .O(N__13498),
            .I(N__13484));
    InMux I__1195 (
            .O(N__13497),
            .I(N__13484));
    InMux I__1194 (
            .O(N__13496),
            .I(N__13484));
    InMux I__1193 (
            .O(N__13495),
            .I(N__13484));
    LocalMux I__1192 (
            .O(N__13484),
            .I(\Inst_eia232.Inst_transmitter.counter_1 ));
    CascadeMux I__1191 (
            .O(N__13481),
            .I(N__13476));
    CascadeMux I__1190 (
            .O(N__13480),
            .I(N__13472));
    InMux I__1189 (
            .O(N__13479),
            .I(N__13465));
    InMux I__1188 (
            .O(N__13476),
            .I(N__13465));
    InMux I__1187 (
            .O(N__13475),
            .I(N__13465));
    InMux I__1186 (
            .O(N__13472),
            .I(N__13462));
    LocalMux I__1185 (
            .O(N__13465),
            .I(\Inst_eia232.Inst_transmitter.counter_2 ));
    LocalMux I__1184 (
            .O(N__13462),
            .I(\Inst_eia232.Inst_transmitter.counter_2 ));
    CEMux I__1183 (
            .O(N__13457),
            .I(N__13454));
    LocalMux I__1182 (
            .O(N__13454),
            .I(N__13451));
    Span4Mux_v I__1181 (
            .O(N__13451),
            .I(N__13448));
    Span4Mux_s0_h I__1180 (
            .O(N__13448),
            .I(N__13445));
    Odrv4 I__1179 (
            .O(N__13445),
            .I(\Inst_eia232.Inst_transmitter.n3594 ));
    CascadeMux I__1178 (
            .O(N__13442),
            .I(\Inst_eia232.Inst_transmitter.n3594_cascade_ ));
    SRMux I__1177 (
            .O(N__13439),
            .I(N__13436));
    LocalMux I__1176 (
            .O(N__13436),
            .I(N__13433));
    Span4Mux_s1_h I__1175 (
            .O(N__13433),
            .I(N__13430));
    Odrv4 I__1174 (
            .O(N__13430),
            .I(\Inst_eia232.Inst_transmitter.n4719 ));
    CEMux I__1173 (
            .O(N__13427),
            .I(N__13423));
    InMux I__1172 (
            .O(N__13426),
            .I(N__13420));
    LocalMux I__1171 (
            .O(N__13423),
            .I(N__13415));
    LocalMux I__1170 (
            .O(N__13420),
            .I(N__13415));
    Odrv4 I__1169 (
            .O(N__13415),
            .I(n3615));
    InMux I__1168 (
            .O(N__13412),
            .I(N__13404));
    InMux I__1167 (
            .O(N__13411),
            .I(N__13401));
    InMux I__1166 (
            .O(N__13410),
            .I(N__13392));
    InMux I__1165 (
            .O(N__13409),
            .I(N__13392));
    InMux I__1164 (
            .O(N__13408),
            .I(N__13392));
    InMux I__1163 (
            .O(N__13407),
            .I(N__13392));
    LocalMux I__1162 (
            .O(N__13404),
            .I(N__13389));
    LocalMux I__1161 (
            .O(N__13401),
            .I(\Inst_eia232.Inst_transmitter.counter_0 ));
    LocalMux I__1160 (
            .O(N__13392),
            .I(\Inst_eia232.Inst_transmitter.counter_0 ));
    Odrv4 I__1159 (
            .O(N__13389),
            .I(\Inst_eia232.Inst_transmitter.counter_0 ));
    CascadeMux I__1158 (
            .O(N__13382),
            .I(n9_cascade_));
    InMux I__1157 (
            .O(N__13379),
            .I(N__13373));
    InMux I__1156 (
            .O(N__13378),
            .I(N__13373));
    LocalMux I__1155 (
            .O(N__13373),
            .I(\Inst_eia232.Inst_transmitter.bits_3 ));
    CascadeMux I__1154 (
            .O(N__13370),
            .I(N__13366));
    CascadeMux I__1153 (
            .O(N__13369),
            .I(N__13362));
    InMux I__1152 (
            .O(N__13366),
            .I(N__13355));
    InMux I__1151 (
            .O(N__13365),
            .I(N__13355));
    InMux I__1150 (
            .O(N__13362),
            .I(N__13355));
    LocalMux I__1149 (
            .O(N__13355),
            .I(\Inst_eia232.Inst_transmitter.bits_2 ));
    InMux I__1148 (
            .O(N__13352),
            .I(N__13349));
    LocalMux I__1147 (
            .O(N__13349),
            .I(n3493));
    CascadeMux I__1146 (
            .O(N__13346),
            .I(n3493_cascade_));
    InMux I__1145 (
            .O(N__13343),
            .I(N__13340));
    LocalMux I__1144 (
            .O(N__13340),
            .I(N__13337));
    Odrv4 I__1143 (
            .O(N__13337),
            .I(n6749));
    InMux I__1142 (
            .O(N__13334),
            .I(N__13327));
    InMux I__1141 (
            .O(N__13333),
            .I(N__13320));
    InMux I__1140 (
            .O(N__13332),
            .I(N__13320));
    InMux I__1139 (
            .O(N__13331),
            .I(N__13320));
    InMux I__1138 (
            .O(N__13330),
            .I(N__13317));
    LocalMux I__1137 (
            .O(N__13327),
            .I(N__13312));
    LocalMux I__1136 (
            .O(N__13320),
            .I(N__13312));
    LocalMux I__1135 (
            .O(N__13317),
            .I(\Inst_eia232.Inst_transmitter.bits_0 ));
    Odrv12 I__1134 (
            .O(N__13312),
            .I(\Inst_eia232.Inst_transmitter.bits_0 ));
    InMux I__1133 (
            .O(N__13307),
            .I(N__13295));
    InMux I__1132 (
            .O(N__13306),
            .I(N__13295));
    InMux I__1131 (
            .O(N__13305),
            .I(N__13295));
    InMux I__1130 (
            .O(N__13304),
            .I(N__13295));
    LocalMux I__1129 (
            .O(N__13295),
            .I(\Inst_eia232.Inst_transmitter.bits_1 ));
    InMux I__1128 (
            .O(N__13292),
            .I(N__13288));
    CEMux I__1127 (
            .O(N__13291),
            .I(N__13285));
    LocalMux I__1126 (
            .O(N__13288),
            .I(N__13282));
    LocalMux I__1125 (
            .O(N__13285),
            .I(n4082));
    Odrv12 I__1124 (
            .O(N__13282),
            .I(n4082));
    CascadeMux I__1123 (
            .O(N__13277),
            .I(n234_cascade_));
    CascadeMux I__1122 (
            .O(N__13274),
            .I(N__13270));
    InMux I__1121 (
            .O(N__13273),
            .I(N__13267));
    InMux I__1120 (
            .O(N__13270),
            .I(N__13264));
    LocalMux I__1119 (
            .O(N__13267),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_9 ));
    LocalMux I__1118 (
            .O(N__13264),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_9 ));
    CascadeMux I__1117 (
            .O(N__13259),
            .I(N__13256));
    InMux I__1116 (
            .O(N__13256),
            .I(N__13253));
    LocalMux I__1115 (
            .O(N__13253),
            .I(n234));
    InMux I__1114 (
            .O(N__13250),
            .I(N__13244));
    InMux I__1113 (
            .O(N__13249),
            .I(N__13244));
    LocalMux I__1112 (
            .O(N__13244),
            .I(byteDone));
    InMux I__1111 (
            .O(N__13241),
            .I(N__13238));
    LocalMux I__1110 (
            .O(N__13238),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_6 ));
    InMux I__1109 (
            .O(N__13235),
            .I(N__13232));
    LocalMux I__1108 (
            .O(N__13232),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_5 ));
    InMux I__1107 (
            .O(N__13229),
            .I(N__13226));
    LocalMux I__1106 (
            .O(N__13226),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_4 ));
    InMux I__1105 (
            .O(N__13223),
            .I(N__13220));
    LocalMux I__1104 (
            .O(N__13220),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_3 ));
    InMux I__1103 (
            .O(N__13217),
            .I(N__13214));
    LocalMux I__1102 (
            .O(N__13214),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_2 ));
    InMux I__1101 (
            .O(N__13211),
            .I(N__13208));
    LocalMux I__1100 (
            .O(N__13208),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_7 ));
    InMux I__1099 (
            .O(N__13205),
            .I(N__13202));
    LocalMux I__1098 (
            .O(N__13202),
            .I(\Inst_eia232.Inst_transmitter.txBuffer_8 ));
    INV \INVInst_core.Inst_sync.synchronizedInput180_i0C  (
            .O(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .I(N__37605));
    INV \INVInst_core.Inst_sync.synchronizedInput180_i4C  (
            .O(\INVInst_core.Inst_sync.synchronizedInput180_i4C_net ),
            .I(N__37594));
    defparam IN_MUX_bfv_6_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_1_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7921 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7906 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7891 ),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7876 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\Inst_core.Inst_sampler.n7955 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\Inst_core.Inst_sampler.n7963 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\Inst_core.Inst_controller.n7852 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\Inst_core.Inst_controller.n7860 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\GENERIC_FIFO_1.n7843 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(\GENERIC_FIFO_1.n7936 ),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\GENERIC_FIFO_1.n7816 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\GENERIC_FIFO_1.n7825 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\GENERIC_FIFO_1.n7944_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\GENERIC_FIFO_1.n7834 ),
            .carryinitout(bfn_1_14_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.paused_91_LC_1_1_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.paused_91_LC_1_1_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.paused_91_LC_1_1_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.paused_91_LC_1_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15482),
            .lcout(\Inst_eia232.Inst_transmitter.paused ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37515),
            .ce(N__15440),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.bits__i0_LC_1_2_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bits__i0_LC_1_2_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.bits__i0_LC_1_2_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.bits__i0_LC_1_2_0  (
            .in0(_gnd_net_),
            .in1(N__13330),
            .in2(_gnd_net_),
            .in3(N__13292),
            .lcout(\Inst_eia232.Inst_transmitter.bits_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37506),
            .ce(),
            .sr(N__16822));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i7_LC_1_3_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i7_LC_1_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i7_LC_1_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i7_LC_1_3_0  (
            .in0(N__14708),
            .in1(N__13211),
            .in2(_gnd_net_),
            .in3(N__16794),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i6_LC_1_3_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i6_LC_1_3_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i6_LC_1_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i6_LC_1_3_1  (
            .in0(N__16791),
            .in1(N__14195),
            .in2(_gnd_net_),
            .in3(N__13241),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i5_LC_1_3_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i5_LC_1_3_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i5_LC_1_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i5_LC_1_3_2  (
            .in0(N__13847),
            .in1(N__13235),
            .in2(_gnd_net_),
            .in3(N__16793),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i4_LC_1_3_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i4_LC_1_3_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i4_LC_1_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i4_LC_1_3_3  (
            .in0(N__16790),
            .in1(N__14015),
            .in2(_gnd_net_),
            .in3(N__13229),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i3_LC_1_3_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i3_LC_1_3_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i3_LC_1_3_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i3_LC_1_3_4  (
            .in0(N__16823),
            .in1(N__13223),
            .in2(_gnd_net_),
            .in3(N__14006),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i2_LC_1_3_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i2_LC_1_3_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i2_LC_1_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i2_LC_1_3_5  (
            .in0(N__16789),
            .in1(N__13898),
            .in2(_gnd_net_),
            .in3(N__13217),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i8_LC_1_3_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i8_LC_1_3_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i8_LC_1_3_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i8_LC_1_3_6  (
            .in0(N__14039),
            .in1(N__13205),
            .in2(_gnd_net_),
            .in3(N__16795),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i9_LC_1_3_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i9_LC_1_3_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i9_LC_1_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i9_LC_1_3_7  (
            .in0(N__16792),
            .in1(N__14474),
            .in2(_gnd_net_),
            .in3(N__13273),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(N__16686),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i1_3_lut_adj_117_LC_1_4_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1_3_lut_adj_117_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1_3_lut_adj_117_LC_1_4_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1_3_lut_adj_117_LC_1_4_0  (
            .in0(N__16249),
            .in1(N__16778),
            .in2(_gnd_net_),
            .in3(N__13249),
            .lcout(n234),
            .ltout(n234_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.state_i1_LC_1_4_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.state_i1_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.state_i1_LC_1_4_1 .LUT_INIT=16'b0100011000000010;
    LogicCell40 \Inst_eia232.Inst_transmitter.state_i1_LC_1_4_1  (
            .in0(N__15983),
            .in1(N__16187),
            .in2(N__13277),
            .in3(N__14089),
            .lcout(state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.writeByte_83_LC_1_4_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.writeByte_83_LC_1_4_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.writeByte_83_LC_1_4_2 .LUT_INIT=16'b0011001100100000;
    LogicCell40 \Inst_eia232.Inst_transmitter.writeByte_83_LC_1_4_2  (
            .in0(N__14090),
            .in1(N__15981),
            .in2(N__16198),
            .in3(N__16783),
            .lcout(writeByte),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i10_LC_1_4_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i10_LC_1_4_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i10_LC_1_4_3 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i10_LC_1_4_3  (
            .in0(N__16779),
            .in1(_gnd_net_),
            .in2(N__13274),
            .in3(N__16717),
            .lcout(\Inst_eia232.Inst_transmitter.txBuffer_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.state_i0_LC_1_4_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.state_i0_LC_1_4_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.state_i0_LC_1_4_4 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \Inst_eia232.Inst_transmitter.state_i0_LC_1_4_4  (
            .in0(N__16031),
            .in1(N__15982),
            .in2(N__13259),
            .in3(N__16191),
            .lcout(state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i28_LC_1_4_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i28_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i28_LC_1_4_5 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i28_LC_1_4_5  (
            .in0(N__15980),
            .in1(N__14225),
            .in2(N__36422),
            .in3(N__21669),
            .lcout(dataBuffer_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i25_LC_1_4_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i25_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i25_LC_1_4_6 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i25_LC_1_4_6  (
            .in0(N__21668),
            .in1(N__36402),
            .in2(N__13994),
            .in3(N__15984),
            .lcout(dataBuffer_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byteDone_81_LC_1_4_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byteDone_81_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byteDone_81_LC_1_4_7 .LUT_INIT=16'b1100101011001111;
    LogicCell40 \Inst_eia232.Inst_transmitter.byteDone_81_LC_1_4_7  (
            .in0(N__13250),
            .in1(N__14108),
            .in2(N__16804),
            .in3(N__13343),
            .lcout(byteDone),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.bytes_i2_LC_1_5_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bytes_i2_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.bytes_i2_LC_1_5_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.bytes_i2_LC_1_5_0  (
            .in0(N__14180),
            .in1(N__14422),
            .in2(_gnd_net_),
            .in3(N__14146),
            .lcout(bytes_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37483),
            .ce(N__13457),
            .sr(N__13439));
    defparam \Inst_eia232.Inst_transmitter.bytes_i0_LC_1_5_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bytes_i0_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.bytes_i0_LC_1_5_1 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \Inst_eia232.Inst_transmitter.bytes_i0_LC_1_5_1  (
            .in0(N__14147),
            .in1(_gnd_net_),
            .in2(N__14423),
            .in3(N__14178),
            .lcout(bytes_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37483),
            .ce(N__13457),
            .sr(N__13439));
    defparam \Inst_eia232.Inst_transmitter.bytes_i1_LC_1_5_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bytes_i1_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.bytes_i1_LC_1_5_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Inst_eia232.Inst_transmitter.bytes_i1_LC_1_5_2  (
            .in0(N__14179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14418),
            .lcout(bytes_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37483),
            .ce(N__13457),
            .sr(N__13439));
    defparam \Inst_eia232.Inst_transmitter.bits__i3_LC_1_6_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bits__i3_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.bits__i3_LC_1_6_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \Inst_eia232.Inst_transmitter.bits__i3_LC_1_6_0  (
            .in0(N__13379),
            .in1(N__13333),
            .in2(N__13370),
            .in3(N__13307),
            .lcout(\Inst_eia232.Inst_transmitter.bits_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(N__13291),
            .sr(N__16815));
    defparam \Inst_eia232.Inst_transmitter.bits__i2_LC_1_6_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bits__i2_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.bits__i2_LC_1_6_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.bits__i2_LC_1_6_1  (
            .in0(N__13306),
            .in1(N__13365),
            .in2(_gnd_net_),
            .in3(N__13334),
            .lcout(\Inst_eia232.Inst_transmitter.bits_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(N__13291),
            .sr(N__16815));
    defparam \Inst_eia232.Inst_transmitter.i2_4_lut_adj_115_LC_1_6_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i2_4_lut_adj_115_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i2_4_lut_adj_115_LC_1_6_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.i2_4_lut_adj_115_LC_1_6_2  (
            .in0(N__13412),
            .in1(N__13530),
            .in2(N__13480),
            .in3(N__13505),
            .lcout(n9),
            .ltout(n9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i936_3_lut_LC_1_6_3.C_ON=1'b0;
    defparam i936_3_lut_LC_1_6_3.SEQ_MODE=4'b0000;
    defparam i936_3_lut_LC_1_6_3.LUT_INIT=16'b1010111110101010;
    LogicCell40 i936_3_lut_LC_1_6_3 (
            .in0(N__16802),
            .in1(_gnd_net_),
            .in2(N__13382),
            .in3(N__13352),
            .lcout(n4082),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i2_4_lut_LC_1_6_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i2_4_lut_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i2_4_lut_LC_1_6_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.i2_4_lut_LC_1_6_4  (
            .in0(N__13378),
            .in1(N__13331),
            .in2(N__13369),
            .in3(N__13304),
            .lcout(n3493),
            .ltout(n3493_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i5585_2_lut_LC_1_6_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i5585_2_lut_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i5585_2_lut_LC_1_6_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i5585_2_lut_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13346),
            .in3(N__16707),
            .lcout(n6749),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.bits__i1_LC_1_6_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bits__i1_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.bits__i1_LC_1_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.bits__i1_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(N__13332),
            .in2(_gnd_net_),
            .in3(N__13305),
            .lcout(\Inst_eia232.Inst_transmitter.bits_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(N__13291),
            .sr(N__16815));
    defparam i1_2_lut_3_lut_LC_1_6_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_1_6_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_1_6_7.LUT_INIT=16'b1110111011111111;
    LogicCell40 i1_2_lut_3_lut_LC_1_6_7 (
            .in0(N__16803),
            .in1(N__18505),
            .in2(_gnd_net_),
            .in3(N__16706),
            .lcout(n3615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.counter__i3_LC_1_7_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.counter__i3_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.counter__i3_LC_1_7_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.counter__i3_LC_1_7_0  (
            .in0(N__13410),
            .in1(N__13532),
            .in2(N__13481),
            .in3(N__13499),
            .lcout(\Inst_eia232.Inst_transmitter.counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37475),
            .ce(N__13427),
            .sr(N__16688));
    defparam \Inst_eia232.Inst_transmitter.i1166_2_lut_LC_1_7_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1166_2_lut_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1166_2_lut_LC_1_7_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1166_2_lut_LC_1_7_1  (
            .in0(N__13496),
            .in1(N__13407),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Inst_eia232.Inst_transmitter.n2201_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.counter__i4_LC_1_7_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.counter__i4_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.counter__i4_LC_1_7_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.counter__i4_LC_1_7_2  (
            .in0(N__13479),
            .in1(N__13531),
            .in2(N__13517),
            .in3(N__13514),
            .lcout(\Inst_eia232.Inst_transmitter.counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37475),
            .ce(N__13427),
            .sr(N__16688));
    defparam \Inst_eia232.Inst_transmitter.counter__i1_LC_1_7_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.counter__i1_LC_1_7_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.counter__i1_LC_1_7_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \Inst_eia232.Inst_transmitter.counter__i1_LC_1_7_3  (
            .in0(N__13497),
            .in1(N__13408),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_eia232.Inst_transmitter.counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37475),
            .ce(N__13427),
            .sr(N__16688));
    defparam \Inst_eia232.Inst_transmitter.i7274_2_lut_LC_1_7_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i7274_2_lut_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i7274_2_lut_LC_1_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i7274_2_lut_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__13495),
            .in2(_gnd_net_),
            .in3(N__13513),
            .lcout(\Inst_eia232.Inst_transmitter.n8642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.counter__i2_LC_1_7_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.counter__i2_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.counter__i2_LC_1_7_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.counter__i2_LC_1_7_5  (
            .in0(N__13498),
            .in1(N__13409),
            .in2(_gnd_net_),
            .in3(N__13475),
            .lcout(\Inst_eia232.Inst_transmitter.counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37475),
            .ce(N__13427),
            .sr(N__16688));
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_4_lut_LC_1_7_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_4_lut_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_4_lut_LC_1_7_6 .LUT_INIT=16'b1111111100110010;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_4_lut_LC_1_7_6  (
            .in0(N__36346),
            .in1(N__15997),
            .in2(N__16070),
            .in3(N__16196),
            .lcout(\Inst_eia232.Inst_transmitter.n3594 ),
            .ltout(\Inst_eia232.Inst_transmitter.n3594_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i3560_2_lut_3_lut_LC_1_7_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i3560_2_lut_3_lut_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i3560_2_lut_3_lut_LC_1_7_7 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i3560_2_lut_3_lut_LC_1_7_7  (
            .in0(N__16197),
            .in1(_gnd_net_),
            .in2(N__13442),
            .in3(N__15998),
            .lcout(\Inst_eia232.Inst_transmitter.n4719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.counter__i0_LC_1_8_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.counter__i0_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.counter__i0_LC_1_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.counter__i0_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__13411),
            .in2(_gnd_net_),
            .in3(N__13426),
            .lcout(\Inst_eia232.Inst_transmitter.counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37474),
            .ce(),
            .sr(N__16687));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i0_LC_1_9_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i0_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i0_LC_1_9_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i0_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__13601),
            .in2(_gnd_net_),
            .in3(N__36399),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37476),
            .ce(N__21682),
            .sr(N__15902));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i4_LC_1_9_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i4_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i4_LC_1_9_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i4_LC_1_9_1  (
            .in0(N__36401),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13589),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37476),
            .ce(N__21682),
            .sr(N__15902));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i5_LC_1_9_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i5_LC_1_9_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i5_LC_1_9_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i5_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__13580),
            .in2(_gnd_net_),
            .in3(N__36400),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37476),
            .ce(N__21682),
            .sr(N__15902));
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i1_LC_1_10_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i1_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.txBuffer_i1_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.txBuffer_i1_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13571),
            .lcout(tx_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37477),
            .ce(N__16685),
            .sr(N__16814));
    defparam \GENERIC_FIFO_1.write_pointer_919__i0_LC_1_11_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i0_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i0_LC_1_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i0_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__16616),
            .in2(_gnd_net_),
            .in3(N__13547),
            .lcout(\GENERIC_FIFO_1.write_pointer_0 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\GENERIC_FIFO_1.n7836 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i1_LC_1_11_1 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i1_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i1_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i1_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__16568),
            .in2(_gnd_net_),
            .in3(N__13544),
            .lcout(\GENERIC_FIFO_1.write_pointer_1 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7836 ),
            .carryout(\GENERIC_FIFO_1.n7837 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i2_LC_1_11_2 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i2_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i2_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i2_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__16516),
            .in2(_gnd_net_),
            .in3(N__13541),
            .lcout(\GENERIC_FIFO_1.write_pointer_2 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7837 ),
            .carryout(\GENERIC_FIFO_1.n7838 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i3_LC_1_11_3 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i3_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i3_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i3_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__16469),
            .in2(_gnd_net_),
            .in3(N__13538),
            .lcout(\GENERIC_FIFO_1.write_pointer_3 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7838 ),
            .carryout(\GENERIC_FIFO_1.n7839 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i4_LC_1_11_4 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i4_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i4_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i4_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__14934),
            .in2(_gnd_net_),
            .in3(N__13535),
            .lcout(\GENERIC_FIFO_1.write_pointer_4 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7839 ),
            .carryout(\GENERIC_FIFO_1.n7840 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i5_LC_1_11_5 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i5_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i5_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i5_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__14863),
            .in2(_gnd_net_),
            .in3(N__13625),
            .lcout(\GENERIC_FIFO_1.write_pointer_5 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7840 ),
            .carryout(\GENERIC_FIFO_1.n7841 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i6_LC_1_11_6 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i6_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i6_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i6_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__17102),
            .in2(_gnd_net_),
            .in3(N__13622),
            .lcout(\GENERIC_FIFO_1.write_pointer_6 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7841 ),
            .carryout(\GENERIC_FIFO_1.n7842 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i7_LC_1_11_7 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i7_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i7_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i7_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__14567),
            .in2(_gnd_net_),
            .in3(N__13619),
            .lcout(\GENERIC_FIFO_1.write_pointer_7 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7842 ),
            .carryout(\GENERIC_FIFO_1.n7843 ),
            .clk(N__37482),
            .ce(N__14981),
            .sr(N__14822));
    defparam \GENERIC_FIFO_1.write_pointer_919__i8_LC_1_12_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.write_pointer_919__i8_LC_1_12_0 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i8_LC_1_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i8_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__14657),
            .in2(_gnd_net_),
            .in3(N__13616),
            .lcout(\GENERIC_FIFO_1.write_pointer_8 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\GENERIC_FIFO_1.n7844 ),
            .clk(N__37489),
            .ce(N__14996),
            .sr(N__14821));
    defparam \GENERIC_FIFO_1.write_pointer_919__i9_LC_1_12_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.write_pointer_919__i9_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.write_pointer_919__i9_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.write_pointer_919__i9_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__14611),
            .in2(_gnd_net_),
            .in3(N__13613),
            .lcout(\GENERIC_FIFO_1.write_pointer_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37489),
            .ce(N__14996),
            .sr(N__14821));
    defparam \GENERIC_FIFO_1.add_6561_2_lut_LC_1_13_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_2_lut_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_2_lut_LC_1_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_2_lut_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__14792),
            .in2(N__13814),
            .in3(_gnd_net_),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_0 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\GENERIC_FIFO_1.n7827 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_3_lut_LC_1_13_1 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_3_lut_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_3_lut_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_3_lut_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__13802),
            .in2(N__14786),
            .in3(N__13610),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_1 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7827 ),
            .carryout(\GENERIC_FIFO_1.n7828 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_4_lut_LC_1_13_2 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_4_lut_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_4_lut_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_4_lut_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__13790),
            .in2(N__15092),
            .in3(N__13607),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_2 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7828 ),
            .carryout(\GENERIC_FIFO_1.n7829 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_5_lut_LC_1_13_3 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_5_lut_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_5_lut_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_5_lut_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__13778),
            .in2(N__15080),
            .in3(N__13604),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_3 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7829 ),
            .carryout(\GENERIC_FIFO_1.n7830 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_6_lut_LC_1_13_4 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_6_lut_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_6_lut_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_6_lut_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__13766),
            .in2(N__15068),
            .in3(N__13700),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_4 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7830 ),
            .carryout(\GENERIC_FIFO_1.n7831 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_7_lut_LC_1_13_5 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_7_lut_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_7_lut_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_7_lut_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__13751),
            .in2(N__15056),
            .in3(N__13697),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_5 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7831 ),
            .carryout(\GENERIC_FIFO_1.n7832 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_8_lut_LC_1_13_6 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_8_lut_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_8_lut_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_8_lut_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__13739),
            .in2(N__15044),
            .in3(N__13694),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_6 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7832 ),
            .carryout(\GENERIC_FIFO_1.n7833 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_9_lut_LC_1_13_7 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_9_lut_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_9_lut_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_9_lut_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__13727),
            .in2(N__15029),
            .in3(N__13691),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_7 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7833 ),
            .carryout(\GENERIC_FIFO_1.n7834 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_10_lut_LC_1_14_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_6561_10_lut_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_10_lut_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_6561_10_lut_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__15017),
            .in2(N__13715),
            .in3(N__13688),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_8 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\GENERIC_FIFO_1.n7835 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_6561_11_lut_LC_1_14_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.add_6561_11_lut_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_6561_11_lut_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \GENERIC_FIFO_1.add_6561_11_lut_LC_1_14_1  (
            .in0(N__13826),
            .in1(N__15005),
            .in2(_gnd_net_),
            .in3(N__13685),
            .lcout(\GENERIC_FIFO_1.level_9_N_876_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i7_4_lut_LC_1_14_2 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i7_4_lut_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i7_4_lut_LC_1_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \GENERIC_FIFO_1.i7_4_lut_LC_1_14_2  (
            .in0(N__13681),
            .in1(N__13667),
            .in2(N__13655),
            .in3(N__13637),
            .lcout(\GENERIC_FIFO_1.n17_adj_1278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i6_1_lut_LC_1_14_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i6_1_lut_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i6_1_lut_LC_1_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i6_1_lut_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14868),
            .lcout(\GENERIC_FIFO_1.n1375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i7282_4_lut_LC_1_14_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i7282_4_lut_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i7282_4_lut_LC_1_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i7282_4_lut_LC_1_14_7  (
            .in0(N__13682),
            .in1(N__13666),
            .in2(N__13654),
            .in3(N__13636),
            .lcout(\GENERIC_FIFO_1.n8650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_2_lut_LC_1_15_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_2_lut_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_2_lut_LC_1_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_2_lut_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__17233),
            .in2(N__16630),
            .in3(_gnd_net_),
            .lcout(\GENERIC_FIFO_1.n12 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\GENERIC_FIFO_1.n7818 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_3_lut_LC_1_15_1 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_3_lut_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_3_lut_LC_1_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_3_lut_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__16575),
            .in2(_gnd_net_),
            .in3(N__13793),
            .lcout(\GENERIC_FIFO_1.n11 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7818 ),
            .carryout(\GENERIC_FIFO_1.n7819 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_4_lut_LC_1_15_2 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_4_lut_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_4_lut_LC_1_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_4_lut_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__16531),
            .in2(_gnd_net_),
            .in3(N__13781),
            .lcout(\GENERIC_FIFO_1.n10 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7819 ),
            .carryout(\GENERIC_FIFO_1.n7820 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_5_lut_LC_1_15_3 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_5_lut_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_5_lut_LC_1_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_5_lut_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__16483),
            .in2(_gnd_net_),
            .in3(N__13769),
            .lcout(\GENERIC_FIFO_1.n9 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7820 ),
            .carryout(\GENERIC_FIFO_1.n7821 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_6_lut_LC_1_15_4 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_6_lut_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_6_lut_LC_1_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_6_lut_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__14938),
            .in2(_gnd_net_),
            .in3(N__13754),
            .lcout(\GENERIC_FIFO_1.n8 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7821 ),
            .carryout(\GENERIC_FIFO_1.n7822 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_7_lut_LC_1_15_5 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_7_lut_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_7_lut_LC_1_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_7_lut_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__14875),
            .in2(_gnd_net_),
            .in3(N__13742),
            .lcout(\GENERIC_FIFO_1.n7 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7822 ),
            .carryout(\GENERIC_FIFO_1.n7823 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_8_lut_LC_1_15_6 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_8_lut_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_8_lut_LC_1_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_8_lut_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__17116),
            .in2(_gnd_net_),
            .in3(N__13730),
            .lcout(\GENERIC_FIFO_1.n6 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7823 ),
            .carryout(\GENERIC_FIFO_1.n7824 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_9_lut_LC_1_15_7 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_9_lut_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_9_lut_LC_1_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_9_lut_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__14572),
            .in2(_gnd_net_),
            .in3(N__13718),
            .lcout(\GENERIC_FIFO_1.n5 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7824 ),
            .carryout(\GENERIC_FIFO_1.n7825 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_10_lut_LC_1_16_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_10_lut_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_10_lut_LC_1_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_10_lut_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__14662),
            .in2(_gnd_net_),
            .in3(N__13703),
            .lcout(\GENERIC_FIFO_1.n4 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\GENERIC_FIFO_1.n7826 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_11_lut_LC_1_16_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_11_lut_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_1_11_lut_LC_1_16_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_1_11_lut_LC_1_16_1  (
            .in0(N__14616),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13829),
            .lcout(\GENERIC_FIFO_1.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i9_1_lut_LC_1_16_2 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i9_1_lut_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i9_1_lut_LC_1_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i9_1_lut_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14661),
            .lcout(\GENERIC_FIFO_1.n1372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i8_1_lut_LC_1_16_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i8_1_lut_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i8_1_lut_LC_1_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i8_1_lut_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14571),
            .lcout(\GENERIC_FIFO_1.n1373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i10_1_lut_LC_1_16_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i10_1_lut_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i10_1_lut_LC_1_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i10_1_lut_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14615),
            .lcout(\GENERIC_FIFO_1.n1371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i8_LC_2_1_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i8_LC_2_1_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i8_LC_2_1_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i8_LC_2_1_0  (
            .in0(_gnd_net_),
            .in1(N__36413),
            .in2(_gnd_net_),
            .in3(N__15999),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37527),
            .ce(N__21655),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i20_3_lut_3_lut_4_lut_LC_2_2_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i20_3_lut_3_lut_4_lut_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i20_3_lut_3_lut_4_lut_LC_2_2_0 .LUT_INIT=16'b1100110000110010;
    LogicCell40 \Inst_eia232.Inst_transmitter.i20_3_lut_3_lut_4_lut_LC_2_2_0  (
            .in0(N__36406),
            .in1(N__15985),
            .in2(N__16069),
            .in3(N__16192),
            .lcout(n4005),
            .ltout(n4005_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i14_LC_2_2_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i14_LC_2_2_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i14_LC_2_2_1 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i14_LC_2_2_1  (
            .in0(N__15986),
            .in1(N__13841),
            .in2(N__13817),
            .in3(N__36410),
            .lcout(dataBuffer_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i22_LC_2_2_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i22_LC_2_2_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i22_LC_2_2_2 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i22_LC_2_2_2  (
            .in0(N__36408),
            .in1(N__13931),
            .in2(N__21657),
            .in3(N__15991),
            .lcout(dataBuffer_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i24_LC_2_2_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i24_LC_2_2_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i24_LC_2_2_3 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i24_LC_2_2_3  (
            .in0(N__15988),
            .in1(N__21611),
            .in2(N__13913),
            .in3(N__36412),
            .lcout(dataBuffer_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i19_LC_2_2_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i19_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i19_LC_2_2_4 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i19_LC_2_2_4  (
            .in0(N__36407),
            .in1(N__13861),
            .in2(N__21656),
            .in3(N__15990),
            .lcout(dataBuffer_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i18_LC_2_2_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i18_LC_2_2_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i18_LC_2_2_5 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i18_LC_2_2_5  (
            .in0(N__15987),
            .in1(N__21610),
            .in2(N__14033),
            .in3(N__36411),
            .lcout(dataBuffer_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.mux_650_i7_3_lut_LC_2_2_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.mux_650_i7_3_lut_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.mux_650_i7_3_lut_LC_2_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.mux_650_i7_3_lut_LC_2_2_6  (
            .in0(N__13921),
            .in1(N__13930),
            .in2(_gnd_net_),
            .in3(N__13960),
            .lcout(\Inst_eia232.Inst_transmitter.n1323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i30_LC_2_2_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i30_LC_2_2_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i30_LC_2_2_7 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i30_LC_2_2_7  (
            .in0(N__15989),
            .in1(N__36409),
            .in2(N__21658),
            .in3(N__13922),
            .lcout(dataBuffer_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byte__i0_LC_2_3_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i0_LC_2_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i0_LC_2_3_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i0_LC_2_3_0  (
            .in0(N__14749),
            .in1(N__13912),
            .in2(N__13964),
            .in3(N__13868),
            .lcout(\Inst_eia232.Inst_transmitter.byte_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(N__14075),
            .sr(N__16232));
    defparam \Inst_eia232.Inst_transmitter.i2444_3_lut_LC_2_3_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i2444_3_lut_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i2444_3_lut_LC_2_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.i2444_3_lut_LC_2_3_1  (
            .in0(N__13889),
            .in1(N__13880),
            .in2(_gnd_net_),
            .in3(N__16128),
            .lcout(\Inst_eia232.Inst_transmitter.n3571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i7532_2_lut_LC_2_3_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i7532_2_lut_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i7532_2_lut_LC_2_3_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i7532_2_lut_LC_2_3_2  (
            .in0(N__16130),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14303),
            .lcout(),
            .ltout(\Inst_eia232.Inst_transmitter.n8854_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byte__i3_LC_2_3_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i3_LC_2_3_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i3_LC_2_3_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i3_LC_2_3_3  (
            .in0(N__13959),
            .in1(N__13862),
            .in2(N__13850),
            .in3(N__14751),
            .lcout(\Inst_eia232.Inst_transmitter.byte_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(N__14075),
            .sr(N__16232));
    defparam \Inst_eia232.Inst_transmitter.i2505_3_lut_LC_2_3_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i2505_3_lut_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i2505_3_lut_LC_2_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i2505_3_lut_LC_2_3_4  (
            .in0(N__16131),
            .in1(N__13840),
            .in2(_gnd_net_),
            .in3(N__14276),
            .lcout(),
            .ltout(\Inst_eia232.Inst_transmitter.n3632_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byte__i6_LC_2_3_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i6_LC_2_3_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i6_LC_2_3_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i6_LC_2_3_5  (
            .in0(_gnd_net_),
            .in1(N__14048),
            .in2(N__14042),
            .in3(N__14752),
            .lcout(\Inst_eia232.Inst_transmitter.byte_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(N__14075),
            .sr(N__16232));
    defparam \Inst_eia232.Inst_transmitter.i7530_2_lut_LC_2_3_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i7530_2_lut_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i7530_2_lut_LC_2_3_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i7530_2_lut_LC_2_3_6  (
            .in0(N__16129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14333),
            .lcout(),
            .ltout(\Inst_eia232.Inst_transmitter.n8851_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byte__i2_LC_2_3_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i2_LC_2_3_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i2_LC_2_3_7 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i2_LC_2_3_7  (
            .in0(N__13958),
            .in1(N__14032),
            .in2(N__14018),
            .in3(N__14750),
            .lcout(\Inst_eia232.Inst_transmitter.byte_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(N__14075),
            .sr(N__16232));
    defparam \Inst_eia232.Inst_transmitter.byte__i1_LC_2_4_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i1_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i1_LC_2_4_0 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i1_LC_2_4_0  (
            .in0(N__13979),
            .in1(N__14753),
            .in2(N__16132),
            .in3(N__14362),
            .lcout(\Inst_eia232.Inst_transmitter.byte_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37498),
            .ce(N__14071),
            .sr(N__16228));
    defparam \Inst_eia232.Inst_transmitter.i3105_2_lut_LC_2_4_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i3105_2_lut_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i3105_2_lut_LC_2_4_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i3105_2_lut_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(N__15951),
            .in2(_gnd_net_),
            .in3(N__16173),
            .lcout(n4248),
            .ltout(n4248_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_130_LC_2_4_2.C_ON=1'b0;
    defparam i1_4_lut_adj_130_LC_2_4_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_130_LC_2_4_2.LUT_INIT=16'b1111000010000000;
    LogicCell40 i1_4_lut_adj_130_LC_2_4_2 (
            .in0(N__14416),
            .in1(N__14144),
            .in2(N__14000),
            .in3(N__14176),
            .lcout(n1336),
            .ltout(n1336_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i5539_2_lut_LC_2_4_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i5539_2_lut_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i5539_2_lut_LC_2_4_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.i5539_2_lut_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13997),
            .in3(N__14059),
            .lcout(\Inst_eia232.Inst_transmitter.n6703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i7569_2_lut_LC_2_4_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i7569_2_lut_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i7569_2_lut_LC_2_4_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i7569_2_lut_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__13990),
            .in2(_gnd_net_),
            .in3(N__13957),
            .lcout(\Inst_eia232.Inst_transmitter.n8847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_2_4_5.C_ON=1'b0;
    defparam i1_4_lut_LC_2_4_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_2_4_5.LUT_INIT=16'b1110000010000000;
    LogicCell40 i1_4_lut_LC_2_4_5 (
            .in0(N__14177),
            .in1(N__14417),
            .in2(N__13973),
            .in3(N__14145),
            .lcout(n1320),
            .ltout(n1320_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i7548_2_lut_LC_2_4_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i7548_2_lut_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i7548_2_lut_LC_2_4_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i7548_2_lut_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14228),
            .in3(N__14224),
            .lcout(),
            .ltout(\Inst_eia232.Inst_transmitter.n8756_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byte__i4_LC_2_4_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i4_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i4_LC_2_4_7 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i4_LC_2_4_7  (
            .in0(N__14754),
            .in1(N__16121),
            .in2(N__14213),
            .in3(N__14210),
            .lcout(\Inst_eia232.Inst_transmitter.byte_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37498),
            .ce(N__14071),
            .sr(N__16228));
    defparam i7565_3_lut_LC_2_5_0.C_ON=1'b0;
    defparam i7565_3_lut_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam i7565_3_lut_LC_2_5_0.LUT_INIT=16'b1111111111011101;
    LogicCell40 i7565_3_lut_LC_2_5_0 (
            .in0(N__14142),
            .in1(N__14412),
            .in2(_gnd_net_),
            .in3(N__14173),
            .lcout(state_1_N_371_1),
            .ltout(state_1_N_371_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i5581_2_lut_LC_2_5_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i5581_2_lut_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i5581_2_lut_LC_2_5_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i5581_2_lut_LC_2_5_1  (
            .in0(N__16178),
            .in1(_gnd_net_),
            .in2(N__14189),
            .in3(_gnd_net_),
            .lcout(\Inst_eia232.Inst_transmitter.n6745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.bytes_2__I_0_i3_3_lut_LC_2_5_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bytes_2__I_0_i3_3_lut_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.bytes_2__I_0_i3_3_lut_LC_2_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.bytes_2__I_0_i3_3_lut_LC_2_5_2  (
            .in0(N__14501),
            .in1(N__14186),
            .in2(_gnd_net_),
            .in3(N__14174),
            .lcout(\Inst_eia232.Inst_transmitter.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.bytes_2__I_0_i1_3_lut_LC_2_5_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.bytes_2__I_0_i1_3_lut_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.bytes_2__I_0_i1_3_lut_LC_2_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.bytes_2__I_0_i1_3_lut_LC_2_5_3  (
            .in0(N__14413),
            .in1(N__14260),
            .in2(_gnd_net_),
            .in3(N__21539),
            .lcout(\Inst_eia232.Inst_transmitter.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i1201_rep_51_2_lut_LC_2_5_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1201_rep_51_2_lut_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1201_rep_51_2_lut_LC_2_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1201_rep_51_2_lut_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(N__14415),
            .in2(_gnd_net_),
            .in3(N__14175),
            .lcout(),
            .ltout(\Inst_eia232.Inst_transmitter.n9218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.disabled_90_LC_2_5_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.disabled_90_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.disabled_90_LC_2_5_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \Inst_eia232.Inst_transmitter.disabled_90_LC_2_5_5  (
            .in0(N__14239),
            .in1(N__14143),
            .in2(N__14117),
            .in3(N__14114),
            .lcout(disabled),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37492),
            .ce(N__14099),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i1_3_lut_LC_2_5_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1_3_lut_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1_3_lut_LC_2_5_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1_3_lut_LC_2_5_6  (
            .in0(N__15967),
            .in1(N__16177),
            .in2(_gnd_net_),
            .in3(N__14088),
            .lcout(\Inst_eia232.Inst_transmitter.n3652 ),
            .ltout(\Inst_eia232.Inst_transmitter.n3652_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i2_3_lut_LC_2_5_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i2_3_lut_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i2_3_lut_LC_2_5_7 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i2_3_lut_LC_2_5_7  (
            .in0(N__14414),
            .in1(_gnd_net_),
            .in2(N__14384),
            .in3(N__14381),
            .lcout(\Inst_eia232.Inst_transmitter.n2580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i1_LC_2_6_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i1_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i1_LC_2_6_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i1_LC_2_6_0  (
            .in0(N__14375),
            .in1(N__21732),
            .in2(N__14363),
            .in3(N__21664),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i2_LC_2_6_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i2_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i2_LC_2_6_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i2_LC_2_6_1  (
            .in0(N__21662),
            .in1(N__14345),
            .in2(N__21742),
            .in3(N__14332),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i3_LC_2_6_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i3_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i3_LC_2_6_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i3_LC_2_6_2  (
            .in0(N__14302),
            .in1(N__21733),
            .in2(N__14318),
            .in3(N__21665),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i6_LC_2_6_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i6_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i6_LC_2_6_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i6_LC_2_6_3  (
            .in0(N__21663),
            .in1(N__14288),
            .in2(N__21743),
            .in3(N__14275),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i1_LC_2_6_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i1_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i1_LC_2_6_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.disabledBuffer_i1_LC_2_6_4  (
            .in0(N__14249),
            .in1(N__21741),
            .in2(N__21676),
            .in3(N__14261),
            .lcout(\Inst_eia232.Inst_transmitter.disabledBuffer_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.disabledGroupsReg_i0_i1_LC_2_6_5 .C_ON=1'b0;
    defparam \Inst_eia232.disabledGroupsReg_i0_i1_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.disabledGroupsReg_i0_i1_LC_2_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.disabledGroupsReg_i0_i1_LC_2_6_5  (
            .in0(N__22291),
            .in1(N__26730),
            .in2(_gnd_net_),
            .in3(N__14248),
            .lcout(disabledGroupsReg_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i3_LC_2_6_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i3_LC_2_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i3_LC_2_6_6 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \Inst_eia232.Inst_transmitter.disabledBuffer_i3_LC_2_6_6  (
            .in0(N__14240),
            .in1(N__21734),
            .in2(N__21677),
            .in3(N__14510),
            .lcout(\Inst_eia232.Inst_transmitter.disabledBuffer_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.disabledGroupsReg_i0_i3_LC_2_6_7 .C_ON=1'b0;
    defparam \Inst_eia232.disabledGroupsReg_i0_i3_LC_2_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.disabledGroupsReg_i0_i3_LC_2_6_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \Inst_eia232.disabledGroupsReg_i0_i3_LC_2_6_7  (
            .in0(N__14509),
            .in1(_gnd_net_),
            .in2(N__22295),
            .in3(N__31398),
            .lcout(disabledGroupsReg_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i2_LC_2_7_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i2_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i2_LC_2_7_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.disabledBuffer_i2_LC_2_7_0  (
            .in0(N__21729),
            .in1(N__14500),
            .in2(N__14486),
            .in3(N__21667),
            .lcout(\Inst_eia232.Inst_transmitter.disabledBuffer_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.disabledGroupsReg_i0_i2_LC_2_7_1 .C_ON=1'b0;
    defparam \Inst_eia232.disabledGroupsReg_i0_i2_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.disabledGroupsReg_i0_i2_LC_2_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.disabledGroupsReg_i0_i2_LC_2_7_1  (
            .in0(N__22277),
            .in1(N__29127),
            .in2(_gnd_net_),
            .in3(N__14482),
            .lcout(disabledGroupsReg_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byte__i7_LC_2_7_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i7_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i7_LC_2_7_3 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i7_LC_2_7_3  (
            .in0(N__14467),
            .in1(N__14758),
            .in2(N__14444),
            .in3(N__16091),
            .lcout(\Inst_eia232.Inst_transmitter.byte_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i5_LC_2_7_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i5_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i5_LC_2_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i5_LC_2_7_4  (
            .in0(N__21889),
            .in1(N__31406),
            .in2(_gnd_net_),
            .in3(N__14773),
            .lcout(maskRegister_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register_80_LC_2_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register_80_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register_80_LC_2_7_5 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register_80_LC_2_7_5  (
            .in0(N__15695),
            .in1(N__14888),
            .in2(_gnd_net_),
            .in3(N__26291),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.match32Register ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_6_i1_1_lut_LC_2_7_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_6_i1_1_lut_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_6_i1_1_lut_LC_2_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_6_i1_1_lut_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17057),
            .lcout(\GENERIC_FIFO_1.level_9_N_925_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i7_LC_2_7_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i7_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.dataBuffer_i7_LC_2_7_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Inst_eia232.Inst_transmitter.dataBuffer_i7_LC_2_7_7  (
            .in0(N__21666),
            .in1(N__14456),
            .in2(N__14443),
            .in3(N__21730),
            .lcout(\Inst_eia232.Inst_transmitter.dataBuffer_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_2_lut_LC_2_8_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_2_lut_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_2_lut_LC_2_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_2_lut_LC_2_8_0  (
            .in0(N__16346),
            .in1(N__17065),
            .in2(_gnd_net_),
            .in3(N__14429),
            .lcout(\GENERIC_FIFO_1.n8779 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\GENERIC_FIFO_1.n7929 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_3_lut_LC_2_8_1 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_3_lut_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_3_lut_LC_2_8_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_3_lut_LC_2_8_1  (
            .in0(N__16343),
            .in1(N__19415),
            .in2(_gnd_net_),
            .in3(N__14426),
            .lcout(\GENERIC_FIFO_1.n8813 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7929 ),
            .carryout(\GENERIC_FIFO_1.n7930 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_4_lut_LC_2_8_2 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_4_lut_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_4_lut_LC_2_8_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_4_lut_LC_2_8_2  (
            .in0(N__16349),
            .in1(N__19343),
            .in2(_gnd_net_),
            .in3(N__14534),
            .lcout(\GENERIC_FIFO_1.n8814 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7930 ),
            .carryout(\GENERIC_FIFO_1.n7931 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_5_lut_LC_2_8_3 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_5_lut_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_5_lut_LC_2_8_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_5_lut_LC_2_8_3  (
            .in0(N__16341),
            .in1(N__18980),
            .in2(_gnd_net_),
            .in3(N__14531),
            .lcout(\GENERIC_FIFO_1.n8815 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7931 ),
            .carryout(\GENERIC_FIFO_1.n7932 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_6_lut_LC_2_8_4 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_6_lut_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_6_lut_LC_2_8_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_6_lut_LC_2_8_4  (
            .in0(N__16347),
            .in1(N__19259),
            .in2(_gnd_net_),
            .in3(N__14528),
            .lcout(\GENERIC_FIFO_1.n8816 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7932 ),
            .carryout(\GENERIC_FIFO_1.n7933 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_7_lut_LC_2_8_5 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_7_lut_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_7_lut_LC_2_8_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_7_lut_LC_2_8_5  (
            .in0(N__16342),
            .in1(N__19190),
            .in2(_gnd_net_),
            .in3(N__14525),
            .lcout(\GENERIC_FIFO_1.n8817 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7933 ),
            .carryout(\GENERIC_FIFO_1.n7934 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_8_lut_LC_2_8_6 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_8_lut_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_8_lut_LC_2_8_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_8_lut_LC_2_8_6  (
            .in0(N__16348),
            .in1(N__19118),
            .in2(_gnd_net_),
            .in3(N__14522),
            .lcout(\GENERIC_FIFO_1.n8818 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7934 ),
            .carryout(\GENERIC_FIFO_1.n7935 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_9_lut_LC_2_8_7 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_9_lut_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_9_lut_LC_2_8_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_9_lut_LC_2_8_7  (
            .in0(N__16340),
            .in1(N__19757),
            .in2(_gnd_net_),
            .in3(N__14519),
            .lcout(\GENERIC_FIFO_1.n8819 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7935 ),
            .carryout(\GENERIC_FIFO_1.n7936 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_10_lut_LC_2_9_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_10_lut_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_10_lut_LC_2_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_10_lut_LC_2_9_0  (
            .in0(N__16345),
            .in1(N__19565),
            .in2(_gnd_net_),
            .in3(N__14516),
            .lcout(\GENERIC_FIFO_1.n8820 ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\GENERIC_FIFO_1.n7937 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_11_lut_LC_2_9_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_11_lut_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_add_4_11_lut_LC_2_9_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_add_4_11_lut_LC_2_9_1  (
            .in0(N__16344),
            .in1(N__17177),
            .in2(_gnd_net_),
            .in3(N__14513),
            .lcout(\GENERIC_FIFO_1.n8821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105_bdd_4_lut_LC_2_9_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105_bdd_4_lut_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105_bdd_4_lut_LC_2_9_2 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.n9105_bdd_4_lut_LC_2_9_2  (
            .in0(N__25500),
            .in1(N__22074),
            .in2(N__28086),
            .in3(N__14810),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3584_1_lut_LC_2_9_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3584_1_lut_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3584_1_lut_LC_2_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3584_1_lut_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14774),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.byte__i5_LC_2_9_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.byte__i5_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.byte__i5_LC_2_9_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \Inst_eia232.Inst_transmitter.byte__i5_LC_2_9_6  (
            .in0(N__14701),
            .in1(N__14759),
            .in2(N__14717),
            .in3(N__16087),
            .lcout(\Inst_eia232.Inst_transmitter.byte_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37480),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i7308_3_lut_LC_2_10_0 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i7308_3_lut_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i7308_3_lut_LC_2_10_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \GENERIC_FIFO_1.i7308_3_lut_LC_2_10_0  (
            .in0(N__16976),
            .in1(N__16925),
            .in2(_gnd_net_),
            .in3(N__17255),
            .lcout(),
            .ltout(\GENERIC_FIFO_1.n8677_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i1_4_lut_LC_2_10_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i1_4_lut_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i1_4_lut_LC_2_10_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \GENERIC_FIFO_1.i1_4_lut_LC_2_10_1  (
            .in0(N__17306),
            .in1(N__16877),
            .in2(N__14690),
            .in3(N__17234),
            .lcout(\GENERIC_FIFO_1.n1396 ),
            .ltout(\GENERIC_FIFO_1.n1396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i2_4_lut_LC_2_10_2 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i2_4_lut_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i2_4_lut_LC_2_10_2 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \GENERIC_FIFO_1.i2_4_lut_LC_2_10_2  (
            .in0(N__36644),
            .in1(N__30154),
            .in2(N__14687),
            .in3(N__15269),
            .lcout(\GENERIC_FIFO_1.fifo_memory_N_983 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i5_LC_2_10_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i5_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i5_LC_2_10_4 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i5_LC_2_10_4  (
            .in0(N__15827),
            .in1(N__20580),
            .in2(N__18695),
            .in3(N__25512),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37484),
            .ce(),
            .sr(N__14684));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i0_LC_2_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i0_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i0_LC_2_11_0 .LUT_INIT=16'b0110010101101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i0_LC_2_11_0  (
            .in0(N__20309),
            .in1(N__20798),
            .in2(N__30357),
            .in3(N__31816),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37491),
            .ce(),
            .sr(N__18791));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_LC_2_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_LC_2_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_LC_2_11_1  (
            .in0(N__22415),
            .in1(N__29789),
            .in2(N__26831),
            .in3(N__14678),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i7_4_lut_adj_122_LC_2_11_2 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i7_4_lut_adj_122_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i7_4_lut_adj_122_LC_2_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i7_4_lut_adj_122_LC_2_11_2  (
            .in0(N__14930),
            .in1(N__14656),
            .in2(N__14617),
            .in3(N__14566),
            .lcout(),
            .ltout(\GENERIC_FIFO_1.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i9_4_lut_LC_2_11_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i9_4_lut_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i9_4_lut_LC_2_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i9_4_lut_LC_2_11_3  (
            .in0(N__17101),
            .in1(N__16468),
            .in2(N__14999),
            .in3(N__14971),
            .lcout(\GENERIC_FIFO_1.n20_adj_1274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i5_1_lut_LC_2_11_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i5_1_lut_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i5_1_lut_LC_2_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i5_1_lut_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14929),
            .lcout(\GENERIC_FIFO_1.n1376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i4_LC_2_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i4_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i4_LC_2_12_0 .LUT_INIT=16'b0001111011010010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i4_LC_2_12_0  (
            .in0(N__28087),
            .in1(N__20598),
            .in2(N__19070),
            .in3(N__15851),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37497),
            .ce(),
            .sr(N__18860));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_adj_70_LC_2_12_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_adj_70_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_adj_70_LC_2_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_adj_70_LC_2_12_1  (
            .in0(N__14903),
            .in1(N__14897),
            .in2(N__16862),
            .in3(N__15212),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i5_2_lut_LC_2_12_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i5_2_lut_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i5_2_lut_LC_2_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \GENERIC_FIFO_1.i5_2_lut_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__16567),
            .in2(_gnd_net_),
            .in3(N__16615),
            .lcout(),
            .ltout(\GENERIC_FIFO_1.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i10_4_lut_LC_2_12_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i10_4_lut_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i10_4_lut_LC_2_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i10_4_lut_LC_2_12_4  (
            .in0(N__14864),
            .in1(N__16517),
            .in2(N__14831),
            .in3(N__14828),
            .lcout(\GENERIC_FIFO_1.n4721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_7715_LC_2_12_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_7715_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_7715_LC_2_12_5 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_7715_LC_2_12_5  (
            .in0(N__23038),
            .in1(N__30432),
            .in2(N__22087),
            .in3(N__22172),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_2_lut_LC_2_13_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_2_lut_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_2_lut_LC_2_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_2_lut_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__14801),
            .in2(N__15239),
            .in3(_gnd_net_),
            .lcout(\GENERIC_FIFO_1.n24 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\GENERIC_FIFO_1.n7809 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_3_lut_LC_2_13_1 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_3_lut_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_3_lut_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_3_lut_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__19466),
            .in2(_gnd_net_),
            .in3(N__14777),
            .lcout(\GENERIC_FIFO_1.n23 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7809 ),
            .carryout(\GENERIC_FIFO_1.n7810 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_4_lut_LC_2_13_2 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_4_lut_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_4_lut_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_4_lut_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__16832),
            .in2(_gnd_net_),
            .in3(N__15083),
            .lcout(\GENERIC_FIFO_1.n22 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7810 ),
            .carryout(\GENERIC_FIFO_1.n7811 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_5_lut_LC_2_13_3 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_5_lut_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_5_lut_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_5_lut_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__19049),
            .in2(_gnd_net_),
            .in3(N__15071),
            .lcout(\GENERIC_FIFO_1.n21 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7811 ),
            .carryout(\GENERIC_FIFO_1.n7812 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_6_lut_LC_2_13_4 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_6_lut_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_6_lut_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_6_lut_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__16841),
            .in2(_gnd_net_),
            .in3(N__15059),
            .lcout(\GENERIC_FIFO_1.n20 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7812 ),
            .carryout(\GENERIC_FIFO_1.n7813 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_7_lut_LC_2_13_5 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_7_lut_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_7_lut_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_7_lut_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__16379),
            .in2(_gnd_net_),
            .in3(N__15047),
            .lcout(\GENERIC_FIFO_1.n19 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7813 ),
            .carryout(\GENERIC_FIFO_1.n7814 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_8_lut_LC_2_13_6 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_8_lut_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_8_lut_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_8_lut_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__19454),
            .in2(_gnd_net_),
            .in3(N__15032),
            .lcout(\GENERIC_FIFO_1.n18_adj_1275 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7814 ),
            .carryout(\GENERIC_FIFO_1.n7815 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_9_lut_LC_2_13_7 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_9_lut_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_9_lut_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_9_lut_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__15218),
            .in2(_gnd_net_),
            .in3(N__15020),
            .lcout(\GENERIC_FIFO_1.n17 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7815 ),
            .carryout(\GENERIC_FIFO_1.n7816 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_10_lut_LC_2_14_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_10_lut_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_10_lut_LC_2_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_10_lut_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__19298),
            .in2(_gnd_net_),
            .in3(N__15011),
            .lcout(\GENERIC_FIFO_1.n16_adj_1273 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\GENERIC_FIFO_1.n7817 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_11_lut_LC_2_14_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_11_lut_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_912_1372_add_1_add_2_11_lut_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_912_1372_add_1_add_2_11_lut_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__17132),
            .in2(_gnd_net_),
            .in3(N__15008),
            .lcout(\GENERIC_FIFO_1.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i7312_4_lut_LC_2_14_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i7312_4_lut_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i7312_4_lut_LC_2_14_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i7312_4_lut_LC_2_14_3  (
            .in0(N__15136),
            .in1(N__15121),
            .in2(N__15230),
            .in3(N__15275),
            .lcout(\GENERIC_FIFO_1.n8681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i1_3_lut_LC_2_14_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i1_3_lut_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i1_3_lut_LC_2_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i1_3_lut_LC_2_14_4  (
            .in0(N__15736),
            .in1(N__17069),
            .in2(_gnd_net_),
            .in3(N__19612),
            .lcout(\GENERIC_FIFO_1.n78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i680_1_lut_LC_2_14_5 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i680_1_lut_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i680_1_lut_LC_2_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.i680_1_lut_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17229),
            .lcout(\GENERIC_FIFO_1.level_9__N_900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i7286_4_lut_LC_2_14_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i7286_4_lut_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i7286_4_lut_LC_2_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i7286_4_lut_LC_2_14_6  (
            .in0(N__15151),
            .in1(N__15163),
            .in2(N__15188),
            .in3(N__15199),
            .lcout(\GENERIC_FIFO_1.n8654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i8_1_lut_LC_2_14_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i8_1_lut_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i8_1_lut_LC_2_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i8_1_lut_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19752),
            .lcout(\GENERIC_FIFO_1.n1418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i6_LC_2_15_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i6_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i6_LC_2_15_0 .LUT_INIT=16'b0101100101101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i6_LC_2_15_0  (
            .in0(N__18758),
            .in1(N__20603),
            .in2(N__15803),
            .in3(N__30461),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37526),
            .ce(),
            .sr(N__18836));
    defparam \GENERIC_FIFO_1.i6_4_lut_LC_2_15_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i6_4_lut_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i6_4_lut_LC_2_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \GENERIC_FIFO_1.i6_4_lut_LC_2_15_1  (
            .in0(N__15203),
            .in1(N__15187),
            .in2(N__15170),
            .in3(N__15152),
            .lcout(),
            .ltout(\GENERIC_FIFO_1.n16_adj_1276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i8_3_lut_LC_2_15_2 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i8_3_lut_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i8_3_lut_LC_2_15_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \GENERIC_FIFO_1.i8_3_lut_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__15140),
            .in2(N__15125),
            .in3(N__15122),
            .lcout(\GENERIC_FIFO_1.n18_adj_1277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i1_4_lut_adj_119_LC_2_15_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i1_4_lut_adj_119_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i1_4_lut_adj_119_LC_2_15_6 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \GENERIC_FIFO_1.i1_4_lut_adj_119_LC_2_15_6  (
            .in0(N__15110),
            .in1(N__36414),
            .in2(N__15104),
            .in3(N__15371),
            .lcout(\GENERIC_FIFO_1.n141 ),
            .ltout(\GENERIC_FIFO_1.n141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i10_3_lut_LC_2_15_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i10_3_lut_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i10_3_lut_LC_2_15_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i10_3_lut_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__17176),
            .in2(N__15365),
            .in3(N__17194),
            .lcout(\GENERIC_FIFO_1.n69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_prescaler.counter_922_923__i2_LC_2_16_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_prescaler.counter_922_923__i2_LC_2_16_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_prescaler.counter_922_923__i2_LC_2_16_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Inst_eia232.Inst_prescaler.counter_922_923__i2_LC_2_16_0  (
            .in0(N__18528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18553),
            .lcout(\Inst_eia232.Inst_prescaler.counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37538),
            .ce(),
            .sr(N__18434));
    defparam \Inst_eia232.Inst_prescaler.counter_922_923__i1_LC_2_16_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_prescaler.counter_922_923__i1_LC_2_16_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_prescaler.counter_922_923__i1_LC_2_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_eia232.Inst_prescaler.counter_922_923__i1_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18527),
            .lcout(\Inst_eia232.Inst_prescaler.counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37538),
            .ce(),
            .sr(N__18434));
    defparam \Inst_eia232.Inst_receiver.bitcount_i2_LC_4_1_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.bitcount_i2_LC_4_1_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.bitcount_i2_LC_4_1_0 .LUT_INIT=16'b1101001011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.bitcount_i2_LC_4_1_0  (
            .in0(N__15293),
            .in1(N__20185),
            .in2(N__15320),
            .in3(N__15337),
            .lcout(\Inst_eia232.Inst_receiver.bitcount_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(N__17717));
    defparam \Inst_eia232.Inst_receiver.i1108_2_lut_3_lut_LC_4_1_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1108_2_lut_3_lut_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1108_2_lut_3_lut_LC_4_1_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \Inst_eia232.Inst_receiver.i1108_2_lut_3_lut_LC_4_1_1  (
            .in0(N__20182),
            .in1(_gnd_net_),
            .in2(N__15338),
            .in3(N__15290),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n2143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.bitcount_i3_LC_4_1_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.bitcount_i3_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.bitcount_i3_LC_4_1_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \Inst_eia232.Inst_receiver.bitcount_i3_LC_4_1_2  (
            .in0(N__15319),
            .in1(_gnd_net_),
            .in2(N__15341),
            .in3(N__15304),
            .lcout(\Inst_eia232.Inst_receiver.bitcount_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(N__17717));
    defparam \Inst_eia232.Inst_receiver.bitcount_i0_LC_4_1_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.bitcount_i0_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.bitcount_i0_LC_4_1_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \Inst_eia232.Inst_receiver.bitcount_i0_LC_4_1_3  (
            .in0(N__20183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15291),
            .lcout(\Inst_eia232.Inst_receiver.bitcount_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(N__17717));
    defparam \Inst_eia232.Inst_receiver.bitcount_i1_LC_4_1_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.bitcount_i1_LC_4_1_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.bitcount_i1_LC_4_1_4 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \Inst_eia232.Inst_receiver.bitcount_i1_LC_4_1_4  (
            .in0(N__15292),
            .in1(N__20184),
            .in2(_gnd_net_),
            .in3(N__15336),
            .lcout(\Inst_eia232.Inst_receiver.bitcount_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(N__17717));
    defparam \Inst_eia232.Inst_receiver.i3_4_lut_adj_79_LC_4_1_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i3_4_lut_adj_79_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i3_4_lut_adj_79_LC_4_1_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \Inst_eia232.Inst_receiver.i3_4_lut_adj_79_LC_4_1_5  (
            .in0(N__15332),
            .in1(N__15315),
            .in2(N__15305),
            .in3(N__15289),
            .lcout(\Inst_eia232.Inst_receiver.n7_adj_1264 ),
            .ltout(\Inst_eia232.Inst_receiver.n7_adj_1264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7493_4_lut_LC_4_1_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7493_4_lut_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7493_4_lut_LC_4_1_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \Inst_eia232.Inst_receiver.i7493_4_lut_LC_4_1_6  (
            .in0(N__15397),
            .in1(N__20181),
            .in2(N__15428),
            .in3(N__15419),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n8769_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i24_4_lut_LC_4_1_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i24_4_lut_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i24_4_lut_LC_4_1_7 .LUT_INIT=16'b1000100000110001;
    LogicCell40 \Inst_eia232.Inst_receiver.i24_4_lut_LC_4_1_7  (
            .in0(N__17861),
            .in1(N__17935),
            .in2(N__15425),
            .in3(N__17674),
            .lcout(n3753),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_4_lut_LC_4_2_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_4_lut_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_4_lut_LC_4_2_0 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_4_lut_LC_4_2_0  (
            .in0(N__20134),
            .in1(N__15511),
            .in2(N__15398),
            .in3(N__15412),
            .lcout(\Inst_eia232.Inst_receiver.n5504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.bytecount_i1_LC_4_2_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.bytecount_i1_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.bytecount_i1_LC_4_2_1 .LUT_INIT=16'b1100110010011100;
    LogicCell40 \Inst_eia232.Inst_receiver.bytecount_i1_LC_4_2_1  (
            .in0(N__20164),
            .in1(N__15395),
            .in2(N__20135),
            .in3(N__20211),
            .lcout(\Inst_eia232.Inst_receiver.bytecount_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37540),
            .ce(N__20098),
            .sr(N__16274));
    defparam \Inst_eia232.Inst_receiver.i5572_2_lut_LC_4_2_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i5572_2_lut_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i5572_2_lut_LC_4_2_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i5572_2_lut_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(N__20129),
            .in2(_gnd_net_),
            .in3(N__20163),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n6736_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.bytecount_i2_LC_4_2_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.bytecount_i2_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.bytecount_i2_LC_4_2_3 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \Inst_eia232.Inst_receiver.bytecount_i2_LC_4_2_3  (
            .in0(N__15413),
            .in1(N__15396),
            .in2(N__15422),
            .in3(N__20212),
            .lcout(\Inst_eia232.Inst_receiver.bytecount_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37540),
            .ce(N__20098),
            .sr(N__16274));
    defparam \Inst_eia232.Inst_receiver.i7495_2_lut_LC_4_2_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7495_2_lut_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7495_2_lut_LC_4_2_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i7495_2_lut_LC_4_2_4  (
            .in0(_gnd_net_),
            .in1(N__20128),
            .in2(_gnd_net_),
            .in3(N__15410),
            .lcout(\Inst_eia232.Inst_receiver.n8772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7214_2_lut_LC_4_2_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7214_2_lut_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7214_2_lut_LC_4_2_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Inst_eia232.Inst_receiver.i7214_2_lut_LC_4_2_5  (
            .in0(N__15411),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15391),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n8582_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7549_4_lut_LC_4_2_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7549_4_lut_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7549_4_lut_LC_4_2_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Inst_eia232.Inst_receiver.i7549_4_lut_LC_4_2_6  (
            .in0(N__20133),
            .in1(N__20209),
            .in2(N__15374),
            .in3(N__20162),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n8831_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i25_4_lut_LC_4_2_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i25_4_lut_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i25_4_lut_LC_4_2_7 .LUT_INIT=16'b1000100001010001;
    LogicCell40 \Inst_eia232.Inst_receiver.i25_4_lut_LC_4_2_7  (
            .in0(N__17976),
            .in1(N__17862),
            .in2(N__15443),
            .in3(N__17673),
            .lcout(\Inst_eia232.Inst_receiver.n3718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i7_LC_4_3_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i7_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i7_LC_4_3_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i7_LC_4_3_0  (
            .in0(N__15509),
            .in1(N__34774),
            .in2(N__15550),
            .in3(N__18228),
            .lcout(cmd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37529),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i6_LC_4_3_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i6_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i6_LC_4_3_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i6_LC_4_3_1  (
            .in0(N__18226),
            .in1(N__15545),
            .in2(N__18375),
            .in3(N__34809),
            .lcout(\Inst_eia232.Inst_receiver.cmd_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37529),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_98_LC_4_3_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_98_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_98_LC_4_3_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_98_LC_4_3_2  (
            .in0(N__15508),
            .in1(N__18364),
            .in2(N__15549),
            .in3(N__18408),
            .lcout(\Inst_eia232.Inst_receiver.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_97_LC_4_3_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_97_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_97_LC_4_3_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_4_lut_adj_97_LC_4_3_3  (
            .in0(N__18363),
            .in1(N__15538),
            .in2(N__18415),
            .in3(N__15506),
            .lcout(\Inst_eia232.Inst_receiver.n14_adj_1265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i8_LC_4_3_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i8_LC_4_3_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i8_LC_4_3_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i8_LC_4_3_4  (
            .in0(N__15510),
            .in1(N__34773),
            .in2(N__18484),
            .in3(N__18229),
            .lcout(nstate_2_N_241_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37529),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_LC_4_3_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_LC_4_3_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_LC_4_3_5  (
            .in0(_gnd_net_),
            .in1(N__15537),
            .in2(_gnd_net_),
            .in3(N__15507),
            .lcout(\Inst_eia232.Inst_receiver.n5498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i4_LC_4_3_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i4_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i4_LC_4_3_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i4_LC_4_3_6  (
            .in0(N__18414),
            .in1(N__18060),
            .in2(N__34839),
            .in3(N__18227),
            .lcout(\Inst_eia232.Inst_receiver.cmd_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37529),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i5_LC_4_3_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i5_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i5_LC_4_3_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i5_LC_4_3_7  (
            .in0(N__18225),
            .in1(N__34805),
            .in2(N__18376),
            .in3(N__18413),
            .lcout(\Inst_eia232.Inst_receiver.cmd_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37529),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_adj_114_LC_4_4_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_adj_114_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_adj_114_LC_4_4_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1_2_lut_adj_114_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__15475),
            .in2(_gnd_net_),
            .in3(N__15452),
            .lcout(\Inst_eia232.Inst_transmitter.n3552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.xon_33_LC_4_4_1 .C_ON=1'b0;
    defparam \Inst_eia232.xon_33_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.xon_33_LC_4_4_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Inst_eia232.xon_33_LC_4_4_1  (
            .in0(N__18310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15461),
            .lcout(\Inst_eia232.xon ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37518),
            .ce(),
            .sr(N__17487));
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i2_LC_4_4_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i2_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i2_LC_4_4_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigcfg__i2_LC_4_4_2  (
            .in0(N__18058),
            .in1(N__18131),
            .in2(N__18203),
            .in3(N__15586),
            .lcout(wrtrigcfg_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37518),
            .ce(),
            .sr(N__17487));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_94_LC_4_4_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_94_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_94_LC_4_4_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_94_LC_4_4_3  (
            .in0(N__18129),
            .in1(N__18193),
            .in2(_gnd_net_),
            .in3(N__18057),
            .lcout(\Inst_eia232.Inst_receiver.n75 ),
            .ltout(\Inst_eia232.Inst_receiver.n75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i2_4_lut_LC_4_4_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i2_4_lut_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i2_4_lut_LC_4_4_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Inst_eia232.Inst_receiver.i2_4_lut_LC_4_4_4  (
            .in0(N__18412),
            .in1(N__18374),
            .in2(N__15464),
            .in3(N__15562),
            .lcout(\Inst_eia232.Inst_receiver.n5597 ),
            .ltout(\Inst_eia232.Inst_receiver.n5597_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.xoff_34_LC_4_4_5 .C_ON=1'b0;
    defparam \Inst_eia232.xoff_34_LC_4_4_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.xoff_34_LC_4_4_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Inst_eia232.xoff_34_LC_4_4_5  (
            .in0(N__18309),
            .in1(_gnd_net_),
            .in2(N__15455),
            .in3(_gnd_net_),
            .lcout(\Inst_eia232.xoff ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37518),
            .ce(),
            .sr(N__17487));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_84_LC_4_4_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_84_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_84_LC_4_4_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_adj_84_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(N__18308),
            .in2(_gnd_net_),
            .in3(N__15631),
            .lcout(\Inst_eia232.Inst_receiver.n90 ),
            .ltout(\Inst_eia232.Inst_receiver.n90_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i1_LC_4_4_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i1_LC_4_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i1_LC_4_4_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigcfg__i1_LC_4_4_7  (
            .in0(N__18130),
            .in1(N__18194),
            .in2(N__15446),
            .in3(N__18059),
            .lcout(wrtrigcfg_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37518),
            .ce(),
            .sr(N__17487));
    defparam \Inst_core.Inst_decoder.wrtrigval__i0_LC_4_5_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigval__i0_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigval__i0_LC_4_5_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigval__i0_LC_4_5_0  (
            .in0(N__15634),
            .in1(N__18295),
            .in2(_gnd_net_),
            .in3(N__17522),
            .lcout(wrtrigval_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(),
            .sr(N__17494));
    defparam \Inst_eia232.id_32_LC_4_5_1 .C_ON=1'b0;
    defparam \Inst_eia232.id_32_LC_4_5_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.id_32_LC_4_5_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Inst_eia232.id_32_LC_4_5_1  (
            .in0(N__18008),
            .in1(N__18339),
            .in2(N__18316),
            .in3(N__15572),
            .lcout(\Inst_eia232.id ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(),
            .sr(N__17494));
    defparam \Inst_core.Inst_decoder.reset_52_LC_4_5_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.reset_52_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.reset_52_LC_4_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Inst_core.Inst_decoder.reset_52_LC_4_5_2  (
            .in0(N__15571),
            .in1(N__18340),
            .in2(N__18017),
            .in3(N__18302),
            .lcout(\Inst_core.resetCmd ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(),
            .sr(N__17494));
    defparam \Inst_core.Inst_decoder.arm_53_LC_4_5_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.arm_53_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.arm_53_LC_4_5_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Inst_core.Inst_decoder.arm_53_LC_4_5_3  (
            .in0(N__17521),
            .in1(N__18338),
            .in2(N__18317),
            .in3(N__15570),
            .lcout(\Inst_core.arm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(),
            .sr(N__17494));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_81_LC_4_5_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_81_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_81_LC_4_5_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_adj_81_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__18293),
            .in2(_gnd_net_),
            .in3(N__18006),
            .lcout(),
            .ltout(n5698_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_decoder.wrFlags_35_LC_4_5_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrFlags_35_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrFlags_35_LC_4_5_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Inst_core.Inst_decoder.wrFlags_35_LC_4_5_5  (
            .in0(N__18341),
            .in1(N__15551),
            .in2(N__15518),
            .in3(N__15515),
            .lcout(wrFlags),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(),
            .sr(N__17494));
    defparam \Inst_core.Inst_decoder.wrtrigmask__i0_LC_4_5_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i0_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i0_LC_4_5_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigmask__i0_LC_4_5_6  (
            .in0(N__15635),
            .in1(N__18294),
            .in2(_gnd_net_),
            .in3(N__18009),
            .lcout(wrtrigmask_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(),
            .sr(N__17494));
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i0_LC_4_5_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i0_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i0_LC_4_5_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigcfg__i0_LC_4_5_7  (
            .in0(N__18007),
            .in1(N__18307),
            .in2(_gnd_net_),
            .in3(N__15633),
            .lcout(wrtrigcfg_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(),
            .sr(N__17494));
    defparam \Inst_core.Inst_decoder.wrtrigval__i2_LC_4_6_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigval__i2_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigval__i2_LC_4_6_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigval__i2_LC_4_6_0  (
            .in0(N__15608),
            .in1(N__18073),
            .in2(N__18200),
            .in3(N__18127),
            .lcout(wrtrigval_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(N__17495));
    defparam \Inst_core.Inst_decoder.wrtrigmask__i3_LC_4_6_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i3_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i3_LC_4_6_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigmask__i3_LC_4_6_1  (
            .in0(N__18126),
            .in1(N__18179),
            .in2(N__18082),
            .in3(N__15604),
            .lcout(wrtrigmask_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(N__17495));
    defparam \Inst_core.Inst_decoder.wrtrigval__i1_LC_4_6_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigval__i1_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigval__i1_LC_4_6_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigval__i1_LC_4_6_2  (
            .in0(N__15605),
            .in1(N__18074),
            .in2(N__18201),
            .in3(N__18122),
            .lcout(wrtrigval_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(N__17495));
    defparam \Inst_core.Inst_decoder.wrtrigmask__i1_LC_4_6_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i1_LC_4_6_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i1_LC_4_6_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigmask__i1_LC_4_6_3  (
            .in0(N__18124),
            .in1(N__18178),
            .in2(N__18081),
            .in3(N__15606),
            .lcout(wrtrigmask_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(N__17495));
    defparam \Inst_core.Inst_decoder.wrtrigmask__i2_LC_4_6_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i2_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigmask__i2_LC_4_6_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigmask__i2_LC_4_6_4  (
            .in0(N__15607),
            .in1(N__18069),
            .in2(N__18199),
            .in3(N__18125),
            .lcout(wrtrigmask_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(N__17495));
    defparam \Inst_eia232.Inst_receiver.i132_2_lut_LC_4_6_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i132_2_lut_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i132_2_lut_LC_4_6_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i132_2_lut_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__18289),
            .in2(_gnd_net_),
            .in3(N__15632),
            .lcout(\Inst_eia232.Inst_receiver.n112 ),
            .ltout(\Inst_eia232.Inst_receiver.n112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_decoder.wrtrigval__i3_LC_4_6_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigval__i3_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigval__i3_LC_4_6_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigval__i3_LC_4_6_6  (
            .in0(N__18177),
            .in1(N__18075),
            .in2(N__15590),
            .in3(N__18128),
            .lcout(wrtrigval_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(N__17495));
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i3_LC_4_6_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i3_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrtrigcfg__i3_LC_4_6_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Inst_core.Inst_decoder.wrtrigcfg__i3_LC_4_6_7  (
            .in0(N__18123),
            .in1(N__15587),
            .in2(N__18083),
            .in3(N__18189),
            .lcout(wrtrigcfg_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(N__17495));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i7_LC_4_7_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i7_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i7_LC_4_7_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i7_LC_4_7_0  (
            .in0(N__34356),
            .in1(N__34820),
            .in2(N__27208),
            .in3(N__34935),
            .lcout(cmd_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37493),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_7_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_7_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i7_LC_4_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i7_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i7_LC_4_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i7_LC_4_7_2  (
            .in0(N__27023),
            .in1(N__27193),
            .in2(_gnd_net_),
            .in3(N__26470),
            .lcout(maskRegister_7_adj_1321),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37493),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i0_LC_4_7_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i0_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i0_LC_4_7_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i0_LC_4_7_3  (
            .in0(N__35956),
            .in1(_gnd_net_),
            .in2(N__20690),
            .in3(N__15718),
            .lcout(valueRegister_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37493),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i31_LC_4_7_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i31_LC_4_7_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i31_LC_4_7_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i31_LC_4_7_4  (
            .in0(N__24049),
            .in1(N__34819),
            .in2(N__20447),
            .in3(N__34934),
            .lcout(cmd_38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37493),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_flags.demux_15_LC_4_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_flags.demux_15_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_flags.demux_15_LC_4_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_flags.demux_15_LC_4_7_5  (
            .in0(N__35955),
            .in1(N__22256),
            .in2(_gnd_net_),
            .in3(N__26244),
            .lcout(flagDemux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37493),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i0_LC_4_7_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i0_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i0_LC_4_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i0_LC_4_7_7  (
            .in0(N__15740),
            .in1(N__17052),
            .in2(_gnd_net_),
            .in3(N__19706),
            .lcout(\GENERIC_FIFO_1.read_pointer_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37493),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i0_LC_4_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i0_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i0_LC_4_8_0 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i0_LC_4_8_0  (
            .in0(N__15872),
            .in1(N__15719),
            .in2(N__20602),
            .in3(N__31796),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37481),
            .ce(),
            .sr(N__20423));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_LC_4_8_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_LC_4_8_1 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister_20__bdd_4_lut_LC_4_8_1  (
            .in0(N__30936),
            .in1(N__32353),
            .in2(N__22088),
            .in3(N__22171),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_bdd_4_lut_LC_4_8_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_bdd_4_lut_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_bdd_4_lut_LC_4_8_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.n9111_bdd_4_lut_LC_4_8_2  (
            .in0(N__33653),
            .in1(N__31795),
            .in2(N__15707),
            .in3(N__22086),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n9114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_762_i1_3_lut_4_lut_LC_4_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_762_i1_3_lut_4_lut_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_762_i1_3_lut_4_lut_LC_4_8_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_762_i1_3_lut_4_lut_LC_4_8_3  (
            .in0(N__21911),
            .in1(N__15668),
            .in2(N__15704),
            .in3(N__24118),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelL16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_LC_4_8_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_LC_4_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3_4_lut_LC_4_8_4  (
            .in0(N__18584),
            .in1(N__20519),
            .in2(N__18614),
            .in3(N__15701),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_706_i1_3_lut_4_lut_LC_4_8_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_706_i1_3_lut_4_lut_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_706_i1_3_lut_4_lut_LC_4_8_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.mux_706_i1_3_lut_4_lut_LC_4_8_5  (
            .in0(N__21910),
            .in1(N__15655),
            .in2(N__15683),
            .in3(N__24119),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.serialChannelH16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i0_LC_4_9_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i0_LC_4_9_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i0_LC_4_9_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i0_LC_4_9_0  (
            .in0(N__26270),
            .in1(N__15667),
            .in2(N__15656),
            .in3(N__18677),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i1_LC_4_9_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i1_LC_4_9_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i1_LC_4_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i1_LC_4_9_1  (
            .in0(N__15651),
            .in1(N__15864),
            .in2(_gnd_net_),
            .in3(N__26263),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i2_LC_4_9_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i2_LC_4_9_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i2_LC_4_9_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i2_LC_4_9_2  (
            .in0(N__26264),
            .in1(_gnd_net_),
            .in2(N__15871),
            .in3(N__20628),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i3_LC_4_9_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i3_LC_4_9_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i3_LC_4_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i3_LC_4_9_3  (
            .in0(N__20629),
            .in1(N__18597),
            .in2(_gnd_net_),
            .in3(N__26265),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i4_LC_4_9_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i4_LC_4_9_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i4_LC_4_9_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i4_LC_4_9_4  (
            .in0(N__26266),
            .in1(_gnd_net_),
            .in2(N__18604),
            .in3(N__18627),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i5_LC_4_9_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i5_LC_4_9_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i5_LC_4_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i5_LC_4_9_5  (
            .in0(N__18628),
            .in1(N__15840),
            .in2(_gnd_net_),
            .in3(N__26267),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i6_LC_4_9_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i6_LC_4_9_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i6_LC_4_9_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i6_LC_4_9_6  (
            .in0(N__26268),
            .in1(_gnd_net_),
            .in2(N__15847),
            .in3(N__15816),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i7_LC_4_9_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i7_LC_4_9_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i7_LC_4_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_i0_i7_LC_4_9_7  (
            .in0(N__15817),
            .in1(N__15793),
            .in2(_gnd_net_),
            .in3(N__26269),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.shiftRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(N__36668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i2_LC_4_10_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i2_LC_4_10_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i2_LC_4_10_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i2_LC_4_10_0  (
            .in0(N__18767),
            .in1(N__22931),
            .in2(_gnd_net_),
            .in3(N__21040),
            .lcout(\Inst_core.Inst_sync.filteredInput_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37501),
            .ce(),
            .sr(N__18716));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i8_3_lut_LC_4_10_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i8_3_lut_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i8_3_lut_LC_4_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i8_3_lut_LC_4_10_1  (
            .in0(N__19774),
            .in1(N__19756),
            .in2(_gnd_net_),
            .in3(N__19704),
            .lcout(\GENERIC_FIFO_1.n71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i9_3_lut_LC_4_10_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i9_3_lut_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i9_3_lut_LC_4_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i9_3_lut_LC_4_10_3  (
            .in0(N__19588),
            .in1(N__19564),
            .in2(_gnd_net_),
            .in3(N__19705),
            .lcout(\GENERIC_FIFO_1.n70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i12_3_lut_LC_4_10_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i12_3_lut_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i12_3_lut_LC_4_10_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Inst_eia232.Inst_receiver.i12_3_lut_LC_4_10_5  (
            .in0(N__17983),
            .in1(N__17884),
            .in2(_gnd_net_),
            .in3(N__17695),
            .lcout(\Inst_eia232.Inst_receiver.n3557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i13_3_lut_LC_4_10_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i13_3_lut_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i13_3_lut_LC_4_10_7 .LUT_INIT=16'b1000100010011001;
    LogicCell40 \Inst_eia232.Inst_receiver.i13_3_lut_LC_4_10_7  (
            .in0(N__17984),
            .in1(N__17885),
            .in2(_gnd_net_),
            .in3(N__17696),
            .lcout(\Inst_eia232.Inst_receiver.n4628 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.busy_87_LC_4_11_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.busy_87_LC_4_11_0 .SEQ_MODE=4'b1001;
    defparam \Inst_eia232.Inst_transmitter.busy_87_LC_4_11_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_eia232.Inst_transmitter.busy_87_LC_4_11_0  (
            .in0(N__16259),
            .in1(N__36425),
            .in2(_gnd_net_),
            .in3(N__16016),
            .lcout(busy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37508),
            .ce(),
            .sr(N__16208));
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_LC_4_11_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_LC_4_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1_2_lut_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__16012),
            .in2(_gnd_net_),
            .in3(N__16206),
            .lcout(\Inst_eia232.Inst_transmitter.n4634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i3103_2_lut_LC_4_11_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i3103_2_lut_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i3103_2_lut_LC_4_11_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i3103_2_lut_LC_4_11_2  (
            .in0(N__16013),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36424),
            .lcout(\Inst_eia232.Inst_transmitter.n4246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_LC_4_11_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_LC_4_11_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i1_2_lut_3_lut_LC_4_11_3  (
            .in0(N__16015),
            .in1(N__16207),
            .in2(_gnd_net_),
            .in3(N__16136),
            .lcout(\Inst_eia232.Inst_transmitter.n8527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i361_2_lut_LC_4_11_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i361_2_lut_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i361_2_lut_LC_4_11_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_eia232.Inst_transmitter.i361_2_lut_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__36423),
            .in2(_gnd_net_),
            .in3(N__16068),
            .lcout(\Inst_eia232.Inst_transmitter.n971 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.i3553_2_lut_LC_4_11_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i3553_2_lut_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i3553_2_lut_LC_4_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.i3553_2_lut_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(N__16014),
            .in2(_gnd_net_),
            .in3(N__21683),
            .lcout(\Inst_eia232.Inst_transmitter.n4712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i2_3_lut_LC_4_11_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i2_3_lut_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i2_3_lut_LC_4_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i2_3_lut_LC_4_11_6  (
            .in0(N__19438),
            .in1(N__19413),
            .in2(_gnd_net_),
            .in3(N__19690),
            .lcout(\GENERIC_FIFO_1.n77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i3_3_lut_LC_4_11_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i3_3_lut_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i3_3_lut_LC_4_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i3_3_lut_LC_4_11_7  (
            .in0(N__19691),
            .in1(N__19360),
            .in2(_gnd_net_),
            .in3(N__19342),
            .lcout(\GENERIC_FIFO_1.n76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i1_LC_4_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i1_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i1_LC_4_12_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i1_LC_4_12_0  (
            .in0(N__22548),
            .in1(N__18773),
            .in2(_gnd_net_),
            .in3(N__22456),
            .lcout(\Inst_core.Inst_sync.filteredInput_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37517),
            .ce(),
            .sr(N__19025));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i4_3_lut_LC_4_12_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i4_3_lut_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i4_3_lut_LC_4_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i4_3_lut_LC_4_12_1  (
            .in0(N__18979),
            .in1(N__19000),
            .in2(_gnd_net_),
            .in3(N__19664),
            .lcout(\GENERIC_FIFO_1.n75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i5_3_lut_LC_4_12_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i5_3_lut_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i5_3_lut_LC_4_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i5_3_lut_LC_4_12_3  (
            .in0(N__19258),
            .in1(N__19282),
            .in2(_gnd_net_),
            .in3(N__19665),
            .lcout(\GENERIC_FIFO_1.n74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i6_3_lut_LC_4_12_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i6_3_lut_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i6_3_lut_LC_4_12_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i6_3_lut_LC_4_12_4  (
            .in0(N__19666),
            .in1(_gnd_net_),
            .in2(N__19186),
            .in3(N__19213),
            .lcout(\GENERIC_FIFO_1.n73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i6_1_lut_LC_4_12_5 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i6_1_lut_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i6_1_lut_LC_4_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i6_1_lut_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19178),
            .lcout(\GENERIC_FIFO_1.n1420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i7_3_lut_LC_4_12_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i7_3_lut_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.read_pointer_921_mux_7_i7_3_lut_LC_4_12_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921_mux_7_i7_3_lut_LC_4_12_6  (
            .in0(N__19667),
            .in1(_gnd_net_),
            .in2(N__19117),
            .in3(N__19135),
            .lcout(\GENERIC_FIFO_1.n72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i6_4_lut_adj_120_LC_4_13_0 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i6_4_lut_adj_120_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i6_4_lut_adj_120_LC_4_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i6_4_lut_adj_120_LC_4_13_0  (
            .in0(N__19182),
            .in1(N__18963),
            .in2(N__19563),
            .in3(N__17056),
            .lcout(),
            .ltout(\GENERIC_FIFO_1.n16_adj_1279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i5619_4_lut_LC_4_13_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i5619_4_lut_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i5619_4_lut_LC_4_13_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \GENERIC_FIFO_1.i5619_4_lut_LC_4_13_1  (
            .in0(N__19248),
            .in1(N__19414),
            .in2(N__16352),
            .in3(N__16847),
            .lcout(\GENERIC_FIFO_1.n142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i7_LC_4_13_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i7_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i7_LC_4_13_2 .LUT_INIT=16'b0001110111100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i7_LC_4_13_2  (
            .in0(N__23037),
            .in1(N__20597),
            .in2(N__16289),
            .in3(N__19040),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37528),
            .ce(),
            .sr(N__18812));
    defparam \GENERIC_FIFO_1.i7_4_lut_adj_121_LC_4_13_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i7_4_lut_adj_121_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i7_4_lut_adj_121_LC_4_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \GENERIC_FIFO_1.i7_4_lut_adj_121_LC_4_13_3  (
            .in0(N__19332),
            .in1(N__19745),
            .in2(N__17172),
            .in3(N__19110),
            .lcout(\GENERIC_FIFO_1.n17_adj_1280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i5_1_lut_LC_4_13_5 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i5_1_lut_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i5_1_lut_LC_4_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i5_1_lut_LC_4_13_5  (
            .in0(N__19247),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\GENERIC_FIFO_1.n1421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i3_1_lut_LC_4_13_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i3_1_lut_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i3_1_lut_LC_4_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i3_1_lut_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19331),
            .lcout(\GENERIC_FIFO_1.n1423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i4_LC_4_14_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i4_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i4_LC_4_14_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i4_LC_4_14_0  (
            .in0(N__21124),
            .in1(N__21151),
            .in2(_gnd_net_),
            .in3(N__19010),
            .lcout(\Inst_core.Inst_sync.filteredInput_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37539),
            .ce(),
            .sr(N__19505));
    defparam \Inst_eia232.Inst_transmitter.i938_2_lut_LC_4_14_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.i938_2_lut_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_transmitter.i938_2_lut_LC_4_14_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Inst_eia232.Inst_transmitter.i938_2_lut_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__16813),
            .in2(_gnd_net_),
            .in3(N__16721),
            .lcout(\Inst_eia232.Inst_transmitter.n3608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.i1047_1_lut_LC_4_14_2 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.i1047_1_lut_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.i1047_1_lut_LC_4_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.i1047_1_lut_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16629),
            .lcout(\GENERIC_FIFO_1.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i2_1_lut_LC_4_14_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i2_1_lut_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i2_1_lut_LC_4_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i2_1_lut_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16579),
            .lcout(\GENERIC_FIFO_1.n1379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i3_1_lut_LC_4_14_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i3_1_lut_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i3_1_lut_LC_4_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i3_1_lut_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16530),
            .lcout(\GENERIC_FIFO_1.n1378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i4_1_lut_LC_4_14_5 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i4_1_lut_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i4_1_lut_LC_4_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i4_1_lut_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16482),
            .lcout(\GENERIC_FIFO_1.n1377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_675_i7_1_lut_LC_4_14_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_675_i7_1_lut_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_675_i7_1_lut_LC_4_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_675_i7_1_lut_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17115),
            .lcout(\GENERIC_FIFO_1.n1374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_2_lut_LC_4_15_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_2_lut_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_2_lut_LC_4_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_676_2_lut_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__17064),
            .in2(N__17018),
            .in3(N__17009),
            .lcout(\GENERIC_FIFO_1.n1391 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\GENERIC_FIFO_1.n7938 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_3_lut_LC_4_15_1 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_3_lut_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_3_lut_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_676_3_lut_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__19390),
            .in2(N__17006),
            .in3(N__16997),
            .lcout(\GENERIC_FIFO_1.n1390 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7938 ),
            .carryout(\GENERIC_FIFO_1.n7939 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_4_lut_LC_4_15_2 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_4_lut_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_4_lut_LC_4_15_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \GENERIC_FIFO_1.add_676_4_lut_LC_4_15_2  (
            .in0(N__16994),
            .in1(N__19319),
            .in2(N__16988),
            .in3(N__16961),
            .lcout(\GENERIC_FIFO_1.n8634 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7939 ),
            .carryout(\GENERIC_FIFO_1.n7940 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_5_lut_LC_4_15_3 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_5_lut_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_5_lut_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_676_5_lut_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__18961),
            .in2(N__16958),
            .in3(N__16949),
            .lcout(\GENERIC_FIFO_1.n1388 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7940 ),
            .carryout(\GENERIC_FIFO_1.n7941 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_6_lut_LC_4_15_4 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_6_lut_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_6_lut_LC_4_15_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \GENERIC_FIFO_1.add_676_6_lut_LC_4_15_4  (
            .in0(N__16946),
            .in1(N__19235),
            .in2(N__16940),
            .in3(N__16910),
            .lcout(\GENERIC_FIFO_1.n8628 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7941 ),
            .carryout(\GENERIC_FIFO_1.n7942 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_7_lut_LC_4_15_5 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_7_lut_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_7_lut_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_676_7_lut_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__16907),
            .in2(N__19177),
            .in3(N__16895),
            .lcout(\GENERIC_FIFO_1.n1386 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7942 ),
            .carryout(\GENERIC_FIFO_1.n7943 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_8_lut_LC_4_15_6 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_8_lut_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_8_lut_LC_4_15_6 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \GENERIC_FIFO_1.add_676_8_lut_LC_4_15_6  (
            .in0(N__16892),
            .in1(N__19098),
            .in2(N__16886),
            .in3(N__16865),
            .lcout(\GENERIC_FIFO_1.n8632 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7943 ),
            .carryout(\GENERIC_FIFO_1.n7944 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_8_THRU_CRY_0_LC_4_15_7 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_8_THRU_CRY_0_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_8_THRU_CRY_0_LC_4_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \GENERIC_FIFO_1.add_676_8_THRU_CRY_0_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__17349),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7944 ),
            .carryout(\GENERIC_FIFO_1.n7944_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_9_lut_LC_4_16_0 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_9_lut_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_9_lut_LC_4_16_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \GENERIC_FIFO_1.add_676_9_lut_LC_4_16_0  (
            .in0(N__17324),
            .in1(N__19729),
            .in2(N__17318),
            .in3(N__17291),
            .lcout(\GENERIC_FIFO_1.n8630 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\GENERIC_FIFO_1.n7945 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_10_lut_LC_4_16_1 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_10_lut_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_10_lut_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \GENERIC_FIFO_1.add_676_10_lut_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__19539),
            .in2(N__17288),
            .in3(N__17276),
            .lcout(\GENERIC_FIFO_1.n1383 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7945 ),
            .carryout(\GENERIC_FIFO_1.n7946 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.add_676_11_lut_LC_4_16_2 .C_ON=1'b1;
    defparam \GENERIC_FIFO_1.add_676_11_lut_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.add_676_11_lut_LC_4_16_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \GENERIC_FIFO_1.add_676_11_lut_LC_4_16_2  (
            .in0(N__17273),
            .in1(N__17152),
            .in2(N__17267),
            .in3(N__17240),
            .lcout(\GENERIC_FIFO_1.n8638 ),
            .ltout(),
            .carryin(\GENERIC_FIFO_1.n7946 ),
            .carryout(\GENERIC_FIFO_1.n1392 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.n1392_THRU_LUT4_0_LC_4_16_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.n1392_THRU_LUT4_0_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.n1392_THRU_LUT4_0_LC_4_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \GENERIC_FIFO_1.n1392_THRU_LUT4_0_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17237),
            .lcout(\GENERIC_FIFO_1.n1392_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i9_LC_4_16_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i9_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i9_LC_4_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i9_LC_4_16_4  (
            .in0(N__19682),
            .in1(N__17201),
            .in2(_gnd_net_),
            .in3(N__17154),
            .lcout(\GENERIC_FIFO_1.read_pointer_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37566),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i10_1_lut_LC_4_16_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i10_1_lut_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i10_1_lut_LC_4_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i10_1_lut_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17153),
            .lcout(\GENERIC_FIFO_1.n1416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_decoder.executePrev_36_LC_5_1_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.executePrev_36_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.executePrev_36_LC_5_1_0 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \Inst_core.Inst_decoder.executePrev_36_LC_5_1_0  (
            .in0(N__17657),
            .in1(_gnd_net_),
            .in2(N__17967),
            .in3(N__17858),
            .lcout(executePrev),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7483_2_lut_LC_5_1_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7483_2_lut_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7483_2_lut_LC_5_1_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Inst_eia232.Inst_receiver.i7483_2_lut_LC_5_1_1  (
            .in0(N__17412),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17653),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n8755_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.state_1__bdd_4_lut_LC_5_1_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.state_1__bdd_4_lut_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.state_1__bdd_4_lut_LC_5_1_2 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \Inst_eia232.Inst_receiver.state_1__bdd_4_lut_LC_5_1_2  (
            .in0(N__17942),
            .in1(N__17856),
            .in2(N__17378),
            .in3(N__17533),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n9123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.state_i1_LC_5_1_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.state_i1_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.state_i1_LC_5_1_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \Inst_eia232.Inst_receiver.state_i1_LC_5_1_3  (
            .in0(N__17860),
            .in1(N__17705),
            .in2(N__17375),
            .in3(N__17366),
            .lcout(\Inst_eia232.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.i5466_2_lut_4_lut_LC_5_1_4 .C_ON=1'b0;
    defparam \Inst_eia232.i5466_2_lut_4_lut_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.i5466_2_lut_4_lut_LC_5_1_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \Inst_eia232.i5466_2_lut_4_lut_LC_5_1_4  (
            .in0(N__17656),
            .in1(N__17372),
            .in2(N__17965),
            .in3(N__17857),
            .lcout(n1917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7487_2_lut_LC_5_1_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7487_2_lut_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7487_2_lut_LC_5_1_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \Inst_eia232.Inst_receiver.i7487_2_lut_LC_5_1_5  (
            .in0(N__17606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17654),
            .lcout(\Inst_eia232.Inst_receiver.n8784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_2_i6_4_lut_LC_5_1_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_2_i6_4_lut_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_2_i6_4_lut_LC_5_1_6 .LUT_INIT=16'b1100010111001111;
    LogicCell40 \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_2_i6_4_lut_LC_5_1_6  (
            .in0(N__17655),
            .in1(N__17534),
            .in2(N__17966),
            .in3(N__17413),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.state_i2_LC_5_1_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.state_i2_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.state_i2_LC_5_1_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \Inst_eia232.Inst_receiver.state_i2_LC_5_1_7  (
            .in0(N__17859),
            .in1(N__17946),
            .in2(N__17360),
            .in3(N__17579),
            .lcout(\Inst_eia232.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i21_3_lut_3_lut_LC_5_2_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i21_3_lut_3_lut_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i21_3_lut_3_lut_LC_5_2_0 .LUT_INIT=16'b0110011001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.i21_3_lut_3_lut_LC_5_2_0  (
            .in0(N__17662),
            .in1(N__17842),
            .in2(_gnd_net_),
            .in3(N__17603),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7647_3_lut_LC_5_2_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7647_3_lut_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7647_3_lut_LC_5_2_1 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \Inst_eia232.Inst_receiver.i7647_3_lut_LC_5_2_1  (
            .in0(N__17937),
            .in1(_gnd_net_),
            .in2(N__17357),
            .in3(N__17395),
            .lcout(\Inst_eia232.Inst_receiver.n4767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i4338_4_lut_LC_5_2_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i4338_4_lut_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i4338_4_lut_LC_5_2_2 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \Inst_eia232.Inst_receiver.i4338_4_lut_LC_5_2_2  (
            .in0(N__20177),
            .in1(N__20210),
            .in2(N__17676),
            .in3(N__17414),
            .lcout(\Inst_eia232.Inst_receiver.n5505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7481_2_lut_3_lut_LC_5_2_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7481_2_lut_3_lut_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7481_2_lut_3_lut_LC_5_2_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \Inst_eia232.Inst_receiver.i7481_2_lut_3_lut_LC_5_2_3  (
            .in0(N__17604),
            .in1(_gnd_net_),
            .in2(N__17863),
            .in3(N__17663),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n8782_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7653_4_lut_LC_5_2_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7653_4_lut_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7653_4_lut_LC_5_2_4 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \Inst_eia232.Inst_receiver.i7653_4_lut_LC_5_2_4  (
            .in0(N__17396),
            .in1(N__18506),
            .in2(N__17399),
            .in3(N__17936),
            .lcout(\Inst_eia232.Inst_receiver.n3676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_adj_99_LC_5_2_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_adj_99_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_adj_99_LC_5_2_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Inst_eia232.Inst_receiver.i2_3_lut_adj_99_LC_5_2_5  (
            .in0(N__17841),
            .in1(N__17661),
            .in2(_gnd_net_),
            .in3(N__20176),
            .lcout(\Inst_eia232.Inst_receiver.n6_adj_1267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_0_i3_4_lut_LC_5_2_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_0_i3_4_lut_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_0_i3_4_lut_LC_5_2_6 .LUT_INIT=16'b1001111100010111;
    LogicCell40 \Inst_eia232.Inst_receiver.state_2__I_0_68_Mux_0_i3_4_lut_LC_5_2_6  (
            .in0(N__17664),
            .in1(N__17938),
            .in2(N__18488),
            .in3(N__17605),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.state_i0_LC_5_2_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.state_i0_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.state_i0_LC_5_2_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \Inst_eia232.Inst_receiver.state_i0_LC_5_2_7  (
            .in0(N__17846),
            .in1(N__17950),
            .in2(N__17387),
            .in3(N__17384),
            .lcout(\Inst_eia232.state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37554),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.counter_925__i3_LC_5_3_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.counter_925__i3_LC_5_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.counter_925__i3_LC_5_3_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.counter_925__i3_LC_5_3_0  (
            .in0(N__17772),
            .in1(N__17744),
            .in2(N__17441),
            .in3(N__17796),
            .lcout(\Inst_eia232.Inst_receiver.counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37542),
            .ce(N__17567),
            .sr(N__17552));
    defparam \Inst_eia232.Inst_receiver.counter_925__i2_LC_5_3_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.counter_925__i2_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.counter_925__i2_LC_5_3_1 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.counter_925__i2_LC_5_3_1  (
            .in0(N__17795),
            .in1(_gnd_net_),
            .in2(N__17747),
            .in3(N__17771),
            .lcout(\Inst_eia232.Inst_receiver.counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37542),
            .ce(N__17567),
            .sr(N__17552));
    defparam \Inst_eia232.Inst_receiver.counter_925__i1_LC_5_3_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.counter_925__i1_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.counter_925__i1_LC_5_3_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Inst_eia232.Inst_receiver.counter_925__i1_LC_5_3_2  (
            .in0(N__17770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17794),
            .lcout(\Inst_eia232.Inst_receiver.counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37542),
            .ce(N__17567),
            .sr(N__17552));
    defparam \Inst_eia232.Inst_receiver.counter_925__i4_LC_5_3_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.counter_925__i4_LC_5_3_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.counter_925__i4_LC_5_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.counter_925__i4_LC_5_3_3  (
            .in0(N__17440),
            .in1(N__17459),
            .in2(_gnd_net_),
            .in3(N__17723),
            .lcout(\Inst_eia232.Inst_receiver.counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37542),
            .ce(N__17567),
            .sr(N__17552));
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_LC_5_3_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_LC_5_3_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \Inst_eia232.Inst_receiver.i2_3_lut_LC_5_3_4  (
            .in0(N__17768),
            .in1(N__17740),
            .in2(_gnd_net_),
            .in3(N__17793),
            .lcout(\Inst_eia232.Inst_receiver.n3504 ),
            .ltout(\Inst_eia232.Inst_receiver.n3504_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_adj_86_LC_5_3_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_adj_86_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i2_3_lut_adj_86_LC_5_3_5 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \Inst_eia232.Inst_receiver.i2_3_lut_adj_86_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(N__17457),
            .in2(N__17570),
            .in3(N__17434),
            .lcout(\Inst_eia232.Inst_receiver.n957 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.counter_925__i0_LC_5_3_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.counter_925__i0_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.counter_925__i0_LC_5_3_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \Inst_eia232.Inst_receiver.counter_925__i0_LC_5_3_6  (
            .in0(N__17769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_eia232.Inst_receiver.counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37542),
            .ce(N__17567),
            .sr(N__17552));
    defparam \Inst_eia232.Inst_receiver.i5570_3_lut_4_lut_LC_5_3_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i5570_3_lut_4_lut_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i5570_3_lut_4_lut_LC_5_3_7 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \Inst_eia232.Inst_receiver.i5570_3_lut_4_lut_LC_5_3_7  (
            .in0(N__17540),
            .in1(N__17458),
            .in2(N__17675),
            .in3(N__17435),
            .lcout(\Inst_eia232.Inst_receiver.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_decoder.wrsize_55_LC_5_4_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrsize_55_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrsize_55_LC_5_4_0 .LUT_INIT=16'b0000001000000010;
    LogicCell40 \Inst_core.Inst_decoder.wrsize_55_LC_5_4_0  (
            .in0(N__17520),
            .in1(N__17503),
            .in2(N__18323),
            .in3(_gnd_net_),
            .lcout(wrsize),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37531),
            .ce(),
            .sr(N__17486));
    defparam \Inst_core.Inst_decoder.wrspeed_54_LC_5_4_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.wrspeed_54_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_decoder.wrspeed_54_LC_5_4_1 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \Inst_core.Inst_decoder.wrspeed_54_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__18319),
            .in2(N__17507),
            .in3(N__18016),
            .lcout(wrDivider),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37531),
            .ce(),
            .sr(N__17486));
    defparam \Inst_core.Inst_sampler.i857_2_lut_LC_5_4_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i857_2_lut_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i857_2_lut_LC_5_4_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_core.Inst_sampler.i857_2_lut_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__30992),
            .in2(_gnd_net_),
            .in3(N__31960),
            .lcout(\Inst_core.Inst_sampler.n1700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i11_4_lut_LC_5_4_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i11_4_lut_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i11_4_lut_LC_5_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i11_4_lut_LC_5_4_3  (
            .in0(N__20269),
            .in1(N__19924),
            .in2(N__20030),
            .in3(N__19975),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.counter_4__I_0_71_i7_2_lut_LC_5_4_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.counter_4__I_0_71_i7_2_lut_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.counter_4__I_0_71_i7_2_lut_LC_5_4_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Inst_eia232.Inst_receiver.counter_4__I_0_71_i7_2_lut_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(N__17456),
            .in2(_gnd_net_),
            .in3(N__17439),
            .lcout(),
            .ltout(\Inst_eia232.Inst_receiver.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i3_4_lut_LC_5_4_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i3_4_lut_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i3_4_lut_LC_5_4_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Inst_eia232.Inst_receiver.i3_4_lut_LC_5_4_5  (
            .in0(N__17797),
            .in1(N__17773),
            .in2(N__17801),
            .in3(N__17745),
            .lcout(\Inst_eia232.Inst_receiver.nstate_2_N_133_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i12_4_lut_LC_5_4_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i12_4_lut_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i12_4_lut_LC_5_4_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i12_4_lut_LC_5_4_6  (
            .in0(N__20251),
            .in1(N__19990),
            .in2(N__20234),
            .in3(N__20284),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i6596_2_lut_3_lut_LC_5_4_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i6596_2_lut_3_lut_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i6596_2_lut_3_lut_LC_5_4_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Inst_eia232.Inst_receiver.i6596_2_lut_3_lut_LC_5_4_7  (
            .in0(N__17798),
            .in1(N__17774),
            .in2(_gnd_net_),
            .in3(N__17746),
            .lcout(\Inst_eia232.Inst_receiver.n7777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i3_LC_5_5_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i3_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i3_LC_5_5_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i3_LC_5_5_0  (
            .in0(N__20507),
            .in1(N__22865),
            .in2(_gnd_net_),
            .in3(N__22435),
            .lcout(\Inst_core.Inst_sync.filteredInput_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37520),
            .ce(),
            .sr(N__18935));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_96_LC_5_5_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_96_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_96_LC_5_5_1 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_96_LC_5_5_1  (
            .in0(N__17694),
            .in1(_gnd_net_),
            .in2(N__17982),
            .in3(N__17882),
            .lcout(\Inst_eia232.Inst_receiver.n3202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i3313_2_lut_LC_5_5_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i3313_2_lut_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i3313_2_lut_LC_5_5_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Inst_eia232.Inst_receiver.i3313_2_lut_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__17971),
            .in2(_gnd_net_),
            .in3(N__17881),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_107_LC_5_5_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_107_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_107_LC_5_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_adj_107_LC_5_5_3  (
            .in0(N__17693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18471),
            .lcout(\Inst_eia232.Inst_receiver.n1_adj_1266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i7571_2_lut_LC_5_5_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i7571_2_lut_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i7571_2_lut_LC_5_5_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i7571_2_lut_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__17692),
            .in2(_gnd_net_),
            .in3(N__17602),
            .lcout(\Inst_eia232.Inst_receiver.n8826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i5549_2_lut_LC_5_5_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i5549_2_lut_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i5549_2_lut_LC_5_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_core.Inst_sampler.i5549_2_lut_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(N__36658),
            .in2(_gnd_net_),
            .in3(N__25367),
            .lcout(\Inst_core.n6713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_prescaler.i5470_2_lut_LC_5_5_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_prescaler.i5470_2_lut_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_prescaler.i5470_2_lut_LC_5_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_eia232.Inst_prescaler.i5470_2_lut_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__18568),
            .in2(_gnd_net_),
            .in3(N__18535),
            .lcout(\Inst_eia232.Inst_prescaler.counter_4__N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_80_LC_5_5_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_80_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_adj_80_LC_5_5_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_adj_80_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(N__18416),
            .in2(_gnd_net_),
            .in3(N__18380),
            .lcout(n12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i3_LC_5_6_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i3_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i3_LC_5_6_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i3_LC_5_6_0  (
            .in0(N__18080),
            .in1(N__18239),
            .in2(N__18202),
            .in3(N__34701),
            .lcout(\Inst_eia232.Inst_receiver.cmd_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i2_LC_5_6_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i2_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i2_LC_5_6_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i2_LC_5_6_1  (
            .in0(N__18237),
            .in1(N__18303),
            .in2(N__18198),
            .in3(N__34706),
            .lcout(\Inst_eia232.Inst_receiver.cmd_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.opcode_i1_LC_5_6_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.opcode_i1_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.opcode_i1_LC_5_6_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.opcode_i1_LC_5_6_2  (
            .in0(N__18114),
            .in1(N__34699),
            .in2(N__18318),
            .in3(N__18238),
            .lcout(\Inst_eia232.Inst_receiver.cmd_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_LC_5_6_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_LC_5_6_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_LC_5_6_3  (
            .in0(N__18173),
            .in1(N__18113),
            .in2(_gnd_net_),
            .in3(N__18079),
            .lcout(\Inst_eia232.Inst_receiver.n69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i27_LC_5_6_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i27_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i27_LC_5_6_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i27_LC_5_6_4  (
            .in0(N__28192),
            .in1(N__35633),
            .in2(N__35067),
            .in3(N__34700),
            .lcout(cmd_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_109_LC_5_6_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_109_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_109_LC_5_6_5 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.i1_2_lut_3_lut_adj_109_LC_5_6_5  (
            .in0(N__17975),
            .in1(N__20091),
            .in2(_gnd_net_),
            .in3(N__17883),
            .lcout(\Inst_eia232.Inst_receiver.n8376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i5_LC_5_6_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i5_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i5_LC_5_6_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i5_LC_5_6_6  (
            .in0(N__29097),
            .in1(N__34698),
            .in2(N__31397),
            .in3(N__35059),
            .lcout(cmd_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_prescaler.scaled_28_LC_5_6_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_prescaler.scaled_28_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_prescaler.scaled_28_LC_5_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_eia232.Inst_prescaler.scaled_28_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__18572),
            .in2(_gnd_net_),
            .in3(N__18539),
            .lcout(trxClock),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i3_LC_5_7_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i3_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i3_LC_5_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i3_LC_5_7_0  (
            .in0(N__26712),
            .in1(N__20689),
            .in2(_gnd_net_),
            .in3(N__18640),
            .lcout(valueRegister_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i3_LC_5_7_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i3_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i3_LC_5_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i3_LC_5_7_1  (
            .in0(N__21865),
            .in1(N__26711),
            .in2(_gnd_net_),
            .in3(N__18895),
            .lcout(maskRegister_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i22_LC_5_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i22_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i22_LC_5_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i22_LC_5_7_2  (
            .in0(N__29757),
            .in1(N__35790),
            .in2(_gnd_net_),
            .in3(N__18735),
            .lcout(configRegister_23_adj_1339),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i22_LC_5_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i22_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i22_LC_5_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i22_LC_5_7_5  (
            .in0(N__26026),
            .in1(N__29758),
            .in2(_gnd_net_),
            .in3(N__18659),
            .lcout(configRegister_23_adj_1379),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i2_LC_5_7_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i2_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i2_LC_5_7_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i2_LC_5_7_6  (
            .in0(N__34817),
            .in1(N__29706),
            .in2(N__34205),
            .in3(N__34996),
            .lcout(cmd_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i32_LC_5_7_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i32_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i32_LC_5_7_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i32_LC_5_7_7  (
            .in0(N__34995),
            .in1(N__20446),
            .in2(N__18470),
            .in3(N__34818),
            .lcout(cmd_39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_7706_LC_5_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_7706_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_7706_LC_5_8_0 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_7706_LC_5_8_0  (
            .in0(N__21818),
            .in1(N__23026),
            .in2(N__30467),
            .in3(N__20410),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_bdd_4_lut_LC_5_8_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_bdd_4_lut_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_bdd_4_lut_LC_5_8_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.n9093_bdd_4_lut_LC_5_8_1  (
            .in0(N__20412),
            .in1(N__28081),
            .in2(N__18437),
            .in3(N__25490),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9096_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_754_i1_3_lut_4_lut_LC_5_8_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_754_i1_3_lut_4_lut_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_754_i1_3_lut_4_lut_LC_5_8_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_754_i1_3_lut_4_lut_LC_5_8_2  (
            .in0(N__21932),
            .in1(N__21466),
            .in2(N__18665),
            .in3(N__18658),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelH16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_LC_5_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_LC_5_8_3 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_20__bdd_4_lut_LC_5_8_3  (
            .in0(N__32343),
            .in1(N__30923),
            .in2(N__20414),
            .in3(N__21817),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_bdd_4_lut_LC_5_8_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_bdd_4_lut_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_bdd_4_lut_LC_5_8_4 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.n9099_bdd_4_lut_LC_5_8_4  (
            .in0(N__33646),
            .in1(N__31794),
            .in2(N__18662),
            .in3(N__20411),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_746_i1_3_lut_4_lut_LC_5_8_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_746_i1_3_lut_4_lut_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_746_i1_3_lut_4_lut_LC_5_8_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.mux_746_i1_3_lut_4_lut_LC_5_8_5  (
            .in0(N__18657),
            .in1(N__21931),
            .in2(N__18644),
            .in3(N__21487),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.serialChannelL16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i3_LC_5_8_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i3_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i3_LC_5_8_6 .LUT_INIT=16'b0110010101101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i3_LC_5_8_6  (
            .in0(N__18641),
            .in1(N__18629),
            .in2(N__20593),
            .in3(N__32344),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37488),
            .ce(),
            .sr(N__18881));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i2_LC_5_9_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i2_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i2_LC_5_9_0 .LUT_INIT=16'b0001110111100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i2_LC_5_9_0  (
            .in0(N__30922),
            .in1(N__20576),
            .in2(N__18605),
            .in3(N__18707),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37504),
            .ce(),
            .sr(N__18911));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_7697_LC_5_9_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_7697_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_7697_LC_5_9_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_7697_LC_5_9_1  (
            .in0(N__20482),
            .in1(N__32338),
            .in2(N__21959),
            .in3(N__30921),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_bdd_4_lut_LC_5_9_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_bdd_4_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_bdd_4_lut_LC_5_9_2 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.n9081_bdd_4_lut_LC_5_9_2  (
            .in0(N__31789),
            .in1(N__33634),
            .in2(N__18578),
            .in3(N__21957),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9084_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_730_i1_3_lut_4_lut_LC_5_9_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_730_i1_3_lut_4_lut_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_730_i1_3_lut_4_lut_LC_5_9_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_730_i1_3_lut_4_lut_LC_5_9_3  (
            .in0(N__18736),
            .in1(N__22108),
            .in2(N__18575),
            .in3(N__24973),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelL16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_LC_5_9_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_LC_5_9_4 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister_20__bdd_4_lut_LC_5_9_4  (
            .in0(N__23025),
            .in1(N__20483),
            .in2(N__30466),
            .in3(N__21956),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_bdd_4_lut_LC_5_9_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_bdd_4_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_bdd_4_lut_LC_5_9_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.n9087_bdd_4_lut_LC_5_9_5  (
            .in0(N__21958),
            .in1(N__28077),
            .in2(N__18740),
            .in3(N__25489),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n9090_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_738_i1_3_lut_4_lut_LC_5_9_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_738_i1_3_lut_4_lut_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_738_i1_3_lut_4_lut_LC_5_9_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.mux_738_i1_3_lut_4_lut_LC_5_9_6  (
            .in0(N__22109),
            .in1(N__18737),
            .in2(N__18719),
            .in3(N__24928),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.serialChannelH16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.i3571_1_lut_LC_5_10_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3571_1_lut_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3571_1_lut_LC_5_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3571_1_lut_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21014),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i0_LC_5_10_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i0_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i0_LC_5_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i0_LC_5_10_1  (
            .in0(N__22025),
            .in1(N__35988),
            .in2(_gnd_net_),
            .in3(N__18800),
            .lcout(maskRegister_0_adj_1288),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i2_LC_5_10_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i2_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i2_LC_5_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i2_LC_5_10_2  (
            .in0(N__20699),
            .in1(N__29714),
            .in2(_gnd_net_),
            .in3(N__18706),
            .lcout(valueRegister_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i23_LC_5_10_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i23_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i23_LC_5_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i23_LC_5_10_3  (
            .in0(N__22226),
            .in1(N__29290),
            .in2(_gnd_net_),
            .in3(N__20845),
            .lcout(configRegister_24_adj_1298),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i24_LC_5_10_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i24_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i24_LC_5_10_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i24_LC_5_10_4  (
            .in0(N__35643),
            .in1(_gnd_net_),
            .in2(N__34098),
            .in3(N__20554),
            .lcout(configRegister_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i5_LC_5_10_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i5_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i5_LC_5_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i5_LC_5_10_5  (
            .in0(N__18691),
            .in1(N__20700),
            .in2(_gnd_net_),
            .in3(N__31369),
            .lcout(valueRegister_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i23_LC_5_10_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i23_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i23_LC_5_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i23_LC_5_10_6  (
            .in0(N__34046),
            .in1(N__18676),
            .in2(_gnd_net_),
            .in3(N__22225),
            .lcout(configRegister_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3483_1_lut_LC_5_10_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3483_1_lut_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3483_1_lut_LC_5_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3483_1_lut_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18799),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i7_LC_5_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i7_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i7_LC_5_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i7_LC_5_11_0  (
            .in0(N__18824),
            .in1(N__27201),
            .in2(_gnd_net_),
            .in3(N__21887),
            .lcout(maskRegister_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i1_LC_5_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i1_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i1_LC_5_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i1_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22558),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i6_LC_5_11_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i6_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i6_LC_5_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i6_LC_5_11_2  (
            .in0(N__34408),
            .in1(N__21886),
            .in2(_gnd_net_),
            .in3(N__18848),
            .lcout(maskRegister_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i2_LC_5_11_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i2_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i2_LC_5_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i2_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22930),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i6_LC_5_11_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i6_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i6_LC_5_11_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i6_LC_5_11_4  (
            .in0(N__34409),
            .in1(N__20695),
            .in2(_gnd_net_),
            .in3(N__18751),
            .lcout(valueRegister_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i7_LC_5_11_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i7_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i7_LC_5_11_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i7_LC_5_11_5  (
            .in0(N__27200),
            .in1(_gnd_net_),
            .in2(N__34501),
            .in3(N__23089),
            .lcout(valueRegister_7_adj_1289),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i2_LC_5_11_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i2_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i2_LC_5_11_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i2_LC_5_11_6  (
            .in0(N__29707),
            .in1(N__21884),
            .in2(_gnd_net_),
            .in3(N__18923),
            .lcout(maskRegister_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i4_LC_5_11_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i4_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i4_LC_5_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i4_LC_5_11_7  (
            .in0(N__21885),
            .in1(N__29110),
            .in2(_gnd_net_),
            .in3(N__18872),
            .lcout(maskRegister_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i0_LC_5_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i0_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i0_LC_5_12_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i0_LC_5_12_0  (
            .in0(N__19514),
            .in1(N__22318),
            .in2(_gnd_net_),
            .in3(N__22636),
            .lcout(\Inst_core.Inst_sync.filteredInput_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37530),
            .ce(),
            .sr(N__20969));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3581_1_lut_LC_5_12_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3581_1_lut_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3581_1_lut_LC_5_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3581_1_lut_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18922),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3582_1_lut_LC_5_12_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3582_1_lut_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3582_1_lut_LC_5_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3582_1_lut_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18896),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3583_1_lut_LC_5_12_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3583_1_lut_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3583_1_lut_LC_5_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3583_1_lut_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18871),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3585_1_lut_LC_5_12_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3585_1_lut_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3585_1_lut_LC_5_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3585_1_lut_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18847),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3586_1_lut_LC_5_12_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3586_1_lut_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3586_1_lut_LC_5_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3586_1_lut_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18823),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_1_lut_LC_5_12_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_1_lut_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_1_lut_LC_5_12_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_1_lut_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__36812),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.n3670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i1_LC_5_13_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i1_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i1_LC_5_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i1_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23302),
            .lcout(\Inst_core.Inst_sync.demuxedInput_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37541),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i7_LC_5_13_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i7_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i7_LC_5_13_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i7_LC_5_13_2  (
            .in0(N__27206),
            .in1(N__22027),
            .in2(_gnd_net_),
            .in3(N__26932),
            .lcout(maskRegister_7_adj_1281),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37541),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i4_LC_5_13_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i4_LC_5_13_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i4_LC_5_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i4_LC_5_13_3  (
            .in0(N__20691),
            .in1(N__19060),
            .in2(_gnd_net_),
            .in3(N__29115),
            .lcout(valueRegister_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37541),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i7_LC_5_13_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i7_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i7_LC_5_13_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i7_LC_5_13_4  (
            .in0(N__27205),
            .in1(N__31111),
            .in2(_gnd_net_),
            .in3(N__24867),
            .lcout(divider_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37541),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i7_LC_5_13_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i7_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i7_LC_5_13_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i7_LC_5_13_5  (
            .in0(N__31110),
            .in1(N__23018),
            .in2(N__22493),
            .in3(N__31964),
            .lcout(memoryOut_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37541),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i2_LC_5_13_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i2_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i2_LC_5_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i2_LC_5_13_6  (
            .in0(N__22026),
            .in1(N__29679),
            .in2(_gnd_net_),
            .in3(N__20909),
            .lcout(maskRegister_2_adj_1286),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37541),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i4_1_lut_LC_5_13_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i4_1_lut_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i4_1_lut_LC_5_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i4_1_lut_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18962),
            .lcout(\GENERIC_FIFO_1.n1422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i7_LC_5_14_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i7_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i7_LC_5_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i7_LC_5_14_0  (
            .in0(N__19036),
            .in1(N__27209),
            .in2(_gnd_net_),
            .in3(N__20701),
            .lcout(valueRegister_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37553),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.i3570_1_lut_LC_5_14_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3570_1_lut_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3570_1_lut_LC_5_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3570_1_lut_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22895),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i4_LC_5_14_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i4_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i4_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i4_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21152),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37553),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i3_LC_5_14_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i3_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i3_LC_5_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i3_LC_5_14_4  (
            .in0(N__19004),
            .in1(N__18969),
            .in2(_gnd_net_),
            .in3(N__19700),
            .lcout(\GENERIC_FIFO_1.read_pointer_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37553),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.i3572_1_lut_LC_5_14_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3572_1_lut_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3572_1_lut_LC_5_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3572_1_lut_LC_5_14_5  (
            .in0(N__22952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i2_1_lut_LC_5_14_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i2_1_lut_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i2_1_lut_LC_5_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i2_1_lut_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19391),
            .lcout(\GENERIC_FIFO_1.n1424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i7_1_lut_LC_5_14_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i7_1_lut_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i7_1_lut_LC_5_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i7_1_lut_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19099),
            .lcout(\GENERIC_FIFO_1.n1419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i1_LC_5_15_0 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i1_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i1_LC_5_15_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i1_LC_5_15_0  (
            .in0(N__19442),
            .in1(N__19400),
            .in2(_gnd_net_),
            .in3(N__19683),
            .lcout(\GENERIC_FIFO_1.read_pointer_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i2_LC_5_15_1 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i2_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i2_LC_5_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i2_LC_5_15_1  (
            .in0(N__19684),
            .in1(N__19364),
            .in2(_gnd_net_),
            .in3(N__19330),
            .lcout(\GENERIC_FIFO_1.read_pointer_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.inv_692_i9_1_lut_LC_5_15_2 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.inv_692_i9_1_lut_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \GENERIC_FIFO_1.inv_692_i9_1_lut_LC_5_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GENERIC_FIFO_1.inv_692_i9_1_lut_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19540),
            .lcout(\GENERIC_FIFO_1.n1417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i4_LC_5_15_3 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i4_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i4_LC_5_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i4_LC_5_15_3  (
            .in0(N__19685),
            .in1(N__19286),
            .in2(_gnd_net_),
            .in3(N__19246),
            .lcout(\GENERIC_FIFO_1.read_pointer_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i5_LC_5_15_4 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i5_LC_5_15_4 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i5_LC_5_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i5_LC_5_15_4  (
            .in0(N__19217),
            .in1(N__19176),
            .in2(_gnd_net_),
            .in3(N__19686),
            .lcout(\GENERIC_FIFO_1.read_pointer_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i6_LC_5_15_5 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i6_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i6_LC_5_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i6_LC_5_15_5  (
            .in0(N__19687),
            .in1(N__19139),
            .in2(_gnd_net_),
            .in3(N__19109),
            .lcout(\GENERIC_FIFO_1.read_pointer_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i7_LC_5_15_6 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i7_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i7_LC_5_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i7_LC_5_15_6  (
            .in0(N__19781),
            .in1(N__19741),
            .in2(_gnd_net_),
            .in3(N__19688),
            .lcout(\GENERIC_FIFO_1.read_pointer_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \GENERIC_FIFO_1.read_pointer_921__i8_LC_5_15_7 .C_ON=1'b0;
    defparam \GENERIC_FIFO_1.read_pointer_921__i8_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \GENERIC_FIFO_1.read_pointer_921__i8_LC_5_15_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \GENERIC_FIFO_1.read_pointer_921__i8_LC_5_15_7  (
            .in0(N__19689),
            .in1(_gnd_net_),
            .in2(N__19553),
            .in3(N__19592),
            .lcout(\GENERIC_FIFO_1.read_pointer_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i0_LC_5_16_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i0_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i0_LC_5_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i0_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22317),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37581),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.i3573_1_lut_LC_5_16_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3573_1_lut_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3573_1_lut_LC_5_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3573_1_lut_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19493),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4732 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i5_LC_5_16_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i5_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i5_LC_5_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input180Delay_i5_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23126),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input180Delay_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37581),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i6_LC_5_16_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i6_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i6_LC_5_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input180Delay_i6_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23165),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input180Delay_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37581),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i4_LC_5_16_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i4_LC_5_16_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i4_LC_5_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i4_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21263),
            .lcout(\Inst_core.Inst_sync.synchronizedInput_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37581),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i4_LC_5_16_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i4_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i4_LC_5_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input180Delay_i4_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21241),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input180Delay_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37581),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i0_LC_5_16_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i0_LC_5_16_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i0_LC_5_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i0_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22685),
            .lcout(\Inst_core.Inst_sync.demuxedInput_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37581),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i1_LC_6_1_0.C_ON=1'b1;
    defparam testcnt_i_917__i1_LC_6_1_0.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i1_LC_6_1_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i1_LC_6_1_0 (
            .in0(_gnd_net_),
            .in1(N__19480),
            .in2(_gnd_net_),
            .in3(N__19469),
            .lcout(testcnt_c_0),
            .ltout(),
            .carryin(bfn_6_1_0_),
            .carryout(n7862),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i2_LC_6_1_1.C_ON=1'b1;
    defparam testcnt_i_917__i2_LC_6_1_1.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i2_LC_6_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i2_LC_6_1_1 (
            .in0(_gnd_net_),
            .in1(N__19903),
            .in2(_gnd_net_),
            .in3(N__19892),
            .lcout(testcnt_c_1),
            .ltout(),
            .carryin(n7862),
            .carryout(n7863),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i3_LC_6_1_2.C_ON=1'b1;
    defparam testcnt_i_917__i3_LC_6_1_2.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i3_LC_6_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i3_LC_6_1_2 (
            .in0(_gnd_net_),
            .in1(N__19882),
            .in2(_gnd_net_),
            .in3(N__19871),
            .lcout(testcnt_c_2),
            .ltout(),
            .carryin(n7863),
            .carryout(n7864),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i4_LC_6_1_3.C_ON=1'b1;
    defparam testcnt_i_917__i4_LC_6_1_3.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i4_LC_6_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i4_LC_6_1_3 (
            .in0(_gnd_net_),
            .in1(N__19867),
            .in2(_gnd_net_),
            .in3(N__19856),
            .lcout(testcnt_c_3),
            .ltout(),
            .carryin(n7864),
            .carryout(n7865),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i5_LC_6_1_4.C_ON=1'b1;
    defparam testcnt_i_917__i5_LC_6_1_4.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i5_LC_6_1_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i5_LC_6_1_4 (
            .in0(_gnd_net_),
            .in1(N__19852),
            .in2(_gnd_net_),
            .in3(N__19841),
            .lcout(testcnt_c_4),
            .ltout(),
            .carryin(n7865),
            .carryout(n7866),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i6_LC_6_1_5.C_ON=1'b1;
    defparam testcnt_i_917__i6_LC_6_1_5.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i6_LC_6_1_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i6_LC_6_1_5 (
            .in0(_gnd_net_),
            .in1(N__19837),
            .in2(_gnd_net_),
            .in3(N__19826),
            .lcout(testcnt_c_5),
            .ltout(),
            .carryin(n7866),
            .carryout(n7867),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i7_LC_6_1_6.C_ON=1'b1;
    defparam testcnt_i_917__i7_LC_6_1_6.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i7_LC_6_1_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i7_LC_6_1_6 (
            .in0(_gnd_net_),
            .in1(N__19816),
            .in2(_gnd_net_),
            .in3(N__19805),
            .lcout(testcnt_c_6),
            .ltout(),
            .carryin(n7867),
            .carryout(n7868),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam testcnt_i_917__i8_LC_6_1_7.C_ON=1'b0;
    defparam testcnt_i_917__i8_LC_6_1_7.SEQ_MODE=4'b1000;
    defparam testcnt_i_917__i8_LC_6_1_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 testcnt_i_917__i8_LC_6_1_7 (
            .in0(_gnd_net_),
            .in1(N__19792),
            .in2(_gnd_net_),
            .in3(N__19802),
            .lcout(testcnt_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i9_LC_6_2_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i9_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i9_LC_6_2_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i9_LC_6_2_0  (
            .in0(N__20011),
            .in1(N__26114),
            .in2(_gnd_net_),
            .in3(N__23998),
            .lcout(configRegister_8_adj_1392),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i2_LC_6_2_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i2_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i2_LC_6_2_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i2_LC_6_2_1  (
            .in0(N__26113),
            .in1(N__19957),
            .in2(_gnd_net_),
            .in3(N__34267),
            .lcout(configRegister_1_adj_1399),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i3_LC_6_2_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i3_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i3_LC_6_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i3_LC_6_2_2  (
            .in0(N__29625),
            .in1(N__19939),
            .in2(_gnd_net_),
            .in3(N__26118),
            .lcout(configRegister_2_adj_1398),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i2_LC_6_2_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i2_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i2_LC_6_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i2_LC_6_2_3  (
            .in0(N__35800),
            .in1(N__23374),
            .in2(_gnd_net_),
            .in3(N__34266),
            .lcout(configRegister_1_adj_1359),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i3_LC_6_2_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i3_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i3_LC_6_2_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i3_LC_6_2_4  (
            .in0(N__29624),
            .in1(N__23344),
            .in2(_gnd_net_),
            .in3(N__35801),
            .lcout(configRegister_2_adj_1358),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i4_LC_6_2_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i4_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i4_LC_6_2_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i4_LC_6_2_5  (
            .in0(N__26721),
            .in1(_gnd_net_),
            .in2(N__26134),
            .in3(N__20053),
            .lcout(configRegister_3_adj_1397),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i4_LC_6_2_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i4_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i4_LC_6_2_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i4_LC_6_2_6  (
            .in0(N__35802),
            .in1(N__23314),
            .in2(_gnd_net_),
            .in3(N__26720),
            .lcout(configRegister_3_adj_1357),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i3_LC_6_2_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i3_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i3_LC_6_2_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i3_LC_6_2_7  (
            .in0(N__29623),
            .in1(N__34776),
            .in2(N__26732),
            .in3(N__35045),
            .lcout(cmd_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i0_LC_6_3_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i0_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i0_LC_6_3_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i0_LC_6_3_0  (
            .in0(N__20498),
            .in1(N__25082),
            .in2(N__21404),
            .in3(N__19961),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_0 ),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7914 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i1_LC_6_3_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i1_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i1_LC_6_3_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i1_LC_6_3_1  (
            .in0(N__19958),
            .in1(N__21437),
            .in2(N__25321),
            .in3(N__19946),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_1 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7914 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7915 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i2_LC_6_3_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i2_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i2_LC_6_3_2 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i2_LC_6_3_2  (
            .in0(N__19943),
            .in1(N__25293),
            .in2(N__19928),
            .in3(N__19913),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_2 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7915 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7916 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i3_LC_6_3_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i3_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i3_LC_6_3_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i3_LC_6_3_3  (
            .in0(N__20054),
            .in1(N__21347),
            .in2(N__25322),
            .in3(N__20042),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_3 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7916 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7917 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i4_LC_6_3_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i4_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i4_LC_6_3_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i4_LC_6_3_4  (
            .in0(N__20465),
            .in1(N__25297),
            .in2(N__21424),
            .in3(N__20039),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_4 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7917 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7918 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i5_LC_6_3_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i5_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i5_LC_6_3_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i5_LC_6_3_5  (
            .in0(N__21287),
            .in1(N__21334),
            .in2(N__25323),
            .in3(N__20036),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_5 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7918 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7919 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i6_LC_6_3_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i6_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i6_LC_6_3_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i6_LC_6_3_6  (
            .in0(N__20354),
            .in1(N__25301),
            .in2(N__21452),
            .in3(N__20033),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_6 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7919 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7920 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i7_LC_6_3_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i7_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i7_LC_6_3_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i7_LC_6_3_7  (
            .in0(N__20324),
            .in1(N__20029),
            .in2(N__25324),
            .in3(N__20015),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_7 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7920 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7921 ),
            .clk(N__37556),
            .ce(N__25697),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i8_LC_6_4_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i8_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i8_LC_6_4_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i8_LC_6_4_0  (
            .in0(N__20012),
            .in1(N__21320),
            .in2(N__25325),
            .in3(N__19997),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_8 ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7922 ),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i9_LC_6_4_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i9_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i9_LC_6_4_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i9_LC_6_4_1  (
            .in0(N__24083),
            .in1(N__25308),
            .in2(N__19994),
            .in3(N__19979),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_9 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7922 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7923 ),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i10_LC_6_4_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i10_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i10_LC_6_4_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i10_LC_6_4_2  (
            .in0(N__21506),
            .in1(N__19976),
            .in2(N__25326),
            .in3(N__19964),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_10 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7923 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7924 ),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i11_LC_6_4_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i11_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i11_LC_6_4_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i11_LC_6_4_3  (
            .in0(N__21518),
            .in1(N__25312),
            .in2(N__20288),
            .in3(N__20273),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_11 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7924 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7925 ),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i12_LC_6_4_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i12_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i12_LC_6_4_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i12_LC_6_4_4  (
            .in0(N__23882),
            .in1(N__20270),
            .in2(N__25327),
            .in3(N__20258),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_12 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7925 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7926 ),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i13_LC_6_4_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i13_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i13_LC_6_4_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i13_LC_6_4_5  (
            .in0(N__26162),
            .in1(N__25316),
            .in2(N__21362),
            .in3(N__20255),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_13 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7926 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7927 ),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i14_LC_6_4_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i14_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i14_LC_6_4_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i14_LC_6_4_6  (
            .in0(N__25547),
            .in1(N__20252),
            .in2(N__25328),
            .in3(N__20240),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_14 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7927 ),
            .carryout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7928 ),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i15_LC_6_4_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i15_LC_6_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i15_LC_6_4_7 .LUT_INIT=16'b1011100001110100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.counter__i15_LC_6_4_7  (
            .in0(N__20233),
            .in1(N__25320),
            .in2(N__21773),
            .in3(N__20237),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37544),
            .ce(N__25696),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.bytecount_i0_LC_6_5_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.bytecount_i0_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.bytecount_i0_LC_6_5_0 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \Inst_eia232.Inst_receiver.bytecount_i0_LC_6_5_0  (
            .in0(N__20115),
            .in1(N__20219),
            .in2(_gnd_net_),
            .in3(N__20186),
            .lcout(\Inst_eia232.Inst_receiver.bytecount_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37533),
            .ce(N__20099),
            .sr(N__20060));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3603_1_lut_LC_6_5_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3603_1_lut_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3603_1_lut_LC_6_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3603_1_lut_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20335),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3604_1_lut_LC_6_5_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3604_1_lut_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3604_1_lut_LC_6_5_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3604_1_lut_LC_6_5_2  (
            .in0(N__20365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3606_1_lut_LC_6_5_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3606_1_lut_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3606_1_lut_LC_6_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3606_1_lut_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20389),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3607_1_lut_LC_6_5_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3607_1_lut_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3607_1_lut_LC_6_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3607_1_lut_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20377),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i6_LC_6_6_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i6_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i6_LC_6_6_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i6_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__34404),
            .in2(N__23921),
            .in3(N__20390),
            .lcout(maskRegister_6_adj_1362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i7_LC_6_6_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i7_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i7_LC_6_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i7_LC_6_6_1  (
            .in0(N__20378),
            .in1(N__27141),
            .in2(_gnd_net_),
            .in3(N__23916),
            .lcout(maskRegister_7_adj_1361),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i4_LC_6_6_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i4_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i4_LC_6_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i4_LC_6_6_2  (
            .in0(N__23912),
            .in1(N__29063),
            .in2(_gnd_net_),
            .in3(N__20366),
            .lcout(maskRegister_4_adj_1364),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i7_LC_6_6_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i7_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i7_LC_6_6_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i7_LC_6_6_3  (
            .in0(N__26048),
            .in1(N__20347),
            .in2(N__34429),
            .in3(_gnd_net_),
            .lcout(configRegister_6_adj_1394),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i3_LC_6_6_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i3_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i3_LC_6_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i3_LC_6_6_4  (
            .in0(N__23911),
            .in1(N__26653),
            .in2(_gnd_net_),
            .in3(N__20336),
            .lcout(maskRegister_3_adj_1365),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i8_LC_6_6_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i8_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i8_LC_6_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i8_LC_6_6_5  (
            .in0(N__26049),
            .in1(N__20320),
            .in2(_gnd_net_),
            .in3(N__27142),
            .lcout(configRegister_7_adj_1393),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i8_LC_6_6_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i8_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i8_LC_6_6_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i8_LC_6_6_6  (
            .in0(N__27140),
            .in1(N__34702),
            .in2(N__23992),
            .in3(N__35058),
            .lcout(cmd_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i9_LC_6_6_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i9_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i9_LC_6_6_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i9_LC_6_6_7  (
            .in0(N__35057),
            .in1(N__23974),
            .in2(N__34777),
            .in3(N__26596),
            .lcout(cmd_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i0_LC_6_7_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i0_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i0_LC_6_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i0_LC_6_7_0  (
            .in0(N__34522),
            .in1(N__35926),
            .in2(_gnd_net_),
            .in3(N__20299),
            .lcout(valueRegister_0_adj_1296),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i3_LC_6_7_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i3_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i3_LC_6_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i3_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22864),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i21_LC_6_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i21_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i21_LC_6_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i21_LC_6_7_2  (
            .in0(N__29331),
            .in1(N__24179),
            .in2(_gnd_net_),
            .in3(N__20721),
            .lcout(configRegister_22_adj_1300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i1_LC_6_7_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i1_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i1_LC_6_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i1_LC_6_7_3  (
            .in0(N__21888),
            .in1(N__34179),
            .in2(_gnd_net_),
            .in3(N__20956),
            .lcout(maskRegister_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i1_LC_6_7_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i1_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i1_LC_6_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i1_LC_6_7_4  (
            .in0(N__26100),
            .in1(N__35927),
            .in2(_gnd_net_),
            .in3(N__20497),
            .lcout(configRegister_0_adj_1400),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i19_LC_6_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i19_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i19_LC_6_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i19_LC_6_7_5  (
            .in0(N__35794),
            .in1(N__26535),
            .in2(_gnd_net_),
            .in3(N__20481),
            .lcout(configRegister_20_adj_1342),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i5_LC_6_7_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i5_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i5_LC_6_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i5_LC_6_7_6  (
            .in0(N__26101),
            .in1(N__20461),
            .in2(_gnd_net_),
            .in3(N__29064),
            .lcout(configRegister_4_adj_1396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i15_LC_6_7_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i15_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i15_LC_6_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i15_LC_6_7_7  (
            .in0(N__35364),
            .in1(N__20445),
            .in2(_gnd_net_),
            .in3(N__22378),
            .lcout(fwd_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3482_1_lut_LC_6_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3482_1_lut_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3482_1_lut_LC_6_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3482_1_lut_LC_6_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21829),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i20_LC_6_8_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i20_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i20_LC_6_8_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i20_LC_6_8_1  (
            .in0(N__24664),
            .in1(N__26119),
            .in2(_gnd_net_),
            .in3(N__20413),
            .lcout(configRegister_21_adj_1381),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i22_LC_6_8_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i22_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i22_LC_6_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i22_LC_6_8_2  (
            .in0(N__29300),
            .in1(N__29751),
            .in2(_gnd_net_),
            .in3(N__20738),
            .lcout(configRegister_23_adj_1299),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i3_LC_6_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i3_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i3_LC_6_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i3_LC_6_8_3  (
            .in0(N__22037),
            .in1(N__26716),
            .in2(_gnd_net_),
            .in3(N__20896),
            .lcout(maskRegister_3_adj_1285),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i20_LC_6_8_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i20_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i20_LC_6_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i20_LC_6_8_4  (
            .in0(N__29299),
            .in1(N__24663),
            .in2(_gnd_net_),
            .in3(N__20763),
            .lcout(configRegister_21_adj_1301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i22_LC_6_8_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i22_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i22_LC_6_8_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i22_LC_6_8_5  (
            .in0(N__24662),
            .in1(N__34775),
            .in2(N__24178),
            .in3(N__34965),
            .lcout(cmd_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i5_LC_6_8_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i5_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i5_LC_6_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i5_LC_6_8_6  (
            .in0(N__34523),
            .in1(N__24328),
            .in2(_gnd_net_),
            .in3(N__31387),
            .lcout(valueRegister_5_adj_1291),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i1_LC_6_8_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i1_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i1_LC_6_8_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.valueRegister_i0_i1_LC_6_8_7  (
            .in0(N__20702),
            .in1(N__34196),
            .in2(_gnd_net_),
            .in3(N__20615),
            .lcout(valueRegister_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_722_i1_3_lut_4_lut_LC_6_9_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_722_i1_3_lut_4_lut_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_722_i1_3_lut_4_lut_LC_6_9_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_722_i1_3_lut_4_lut_LC_6_9_0  (
            .in0(N__20737),
            .in1(N__20774),
            .in2(N__20819),
            .in3(N__20723),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelH16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i1_LC_6_9_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i1_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i1_LC_6_9_1 .LUT_INIT=16'b0110011000111100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_i1_LC_6_9_1  (
            .in0(N__20633),
            .in1(N__20614),
            .in2(N__33652),
            .in3(N__20561),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.intermediateRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37513),
            .ce(),
            .sr(N__20942));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_LC_6_9_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_LC_6_9_2 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_LC_6_9_2  (
            .in0(N__23039),
            .in1(N__20863),
            .in2(N__20765),
            .in3(N__30456),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_bdd_4_lut_LC_6_9_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_bdd_4_lut_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_bdd_4_lut_LC_6_9_3 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.n9075_bdd_4_lut_LC_6_9_3  (
            .in0(N__25488),
            .in1(N__28028),
            .in2(N__20777),
            .in3(N__20762),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_7688_LC_6_9_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_7688_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_7688_LC_6_9_4 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister_20__bdd_4_lut_7688_LC_6_9_4  (
            .in0(N__30924),
            .in1(N__32339),
            .in2(N__20764),
            .in3(N__20862),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_bdd_4_lut_LC_6_9_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_bdd_4_lut_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_bdd_4_lut_LC_6_9_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.n9069_bdd_4_lut_LC_6_9_5  (
            .in0(N__31790),
            .in1(N__33638),
            .in2(N__20768),
            .in3(N__20761),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_714_i1_3_lut_4_lut_LC_6_9_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_714_i1_3_lut_4_lut_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_714_i1_3_lut_4_lut_LC_6_9_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.mux_714_i1_3_lut_4_lut_LC_6_9_6  (
            .in0(N__20736),
            .in1(N__20722),
            .in2(N__20705),
            .in3(N__20833),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.serialChannelL16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_flags.filter_16_LC_6_10_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_flags.filter_16_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_flags.filter_16_LC_6_10_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_flags.filter_16_LC_6_10_0  (
            .in0(N__34226),
            .in1(N__22260),
            .in2(_gnd_net_),
            .in3(N__22583),
            .lcout(flagFilter),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i5_LC_6_10_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i5_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i5_LC_6_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i5_LC_6_10_1  (
            .in0(N__22035),
            .in1(N__31368),
            .in2(_gnd_net_),
            .in3(N__20878),
            .lcout(maskRegister_5_adj_1283),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i4_LC_6_10_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i4_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i4_LC_6_10_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i4_LC_6_10_2  (
            .in0(N__35365),
            .in1(N__26519),
            .in2(N__24239),
            .in3(_gnd_net_),
            .lcout(fwd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i4_LC_6_10_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i4_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i4_LC_6_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i4_LC_6_10_3  (
            .in0(N__29109),
            .in1(N__34529),
            .in2(_gnd_net_),
            .in3(N__24550),
            .lcout(valueRegister_4_adj_1292),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i1_LC_6_10_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i1_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i1_LC_6_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i1_LC_6_10_4  (
            .in0(N__34227),
            .in1(N__22034),
            .in2(_gnd_net_),
            .in3(N__20923),
            .lcout(maskRegister_1_adj_1287),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i21_LC_6_10_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i21_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i21_LC_6_10_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i21_LC_6_10_5  (
            .in0(N__26518),
            .in1(N__34841),
            .in2(N__24684),
            .in3(N__35056),
            .lcout(cmd_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i23_LC_6_10_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i23_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i23_LC_6_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i23_LC_6_10_6  (
            .in0(N__35832),
            .in1(N__24949),
            .in2(_gnd_net_),
            .in3(N__22218),
            .lcout(configRegister_24_adj_1338),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i19_LC_6_10_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i19_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i19_LC_6_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i19_LC_6_10_7  (
            .in0(N__26520),
            .in1(N__29326),
            .in2(_gnd_net_),
            .in3(N__20864),
            .lcout(configRegister_20_adj_1302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i0_LC_6_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i0_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i0_LC_6_11_0 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i0_LC_6_11_0  (
            .in0(N__26356),
            .in1(N__20818),
            .in2(N__20849),
            .in3(N__20834),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i1_LC_6_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i1_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i1_LC_6_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i1_LC_6_11_1  (
            .in0(N__20817),
            .in1(N__20790),
            .in2(_gnd_net_),
            .in3(N__26349),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i2_LC_6_11_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i2_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i2_LC_6_11_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i2_LC_6_11_2  (
            .in0(N__26350),
            .in1(_gnd_net_),
            .in2(N__20797),
            .in3(N__22122),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i3_LC_6_11_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i3_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i3_LC_6_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i3_LC_6_11_3  (
            .in0(N__22123),
            .in1(N__29802),
            .in2(_gnd_net_),
            .in3(N__26351),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i4_LC_6_11_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i4_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i4_LC_6_11_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i4_LC_6_11_4  (
            .in0(N__26352),
            .in1(_gnd_net_),
            .in2(N__29809),
            .in3(N__26856),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i5_LC_6_11_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i5_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i5_LC_6_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i5_LC_6_11_5  (
            .in0(N__26857),
            .in1(N__24573),
            .in2(_gnd_net_),
            .in3(N__26353),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i6_LC_6_11_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i6_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i6_LC_6_11_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i6_LC_6_11_6  (
            .in0(N__26354),
            .in1(_gnd_net_),
            .in2(N__24580),
            .in3(N__24309),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i7_LC_6_11_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i7_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i7_LC_6_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_i0_i7_LC_6_11_7  (
            .in0(N__24310),
            .in1(N__30244),
            .in2(_gnd_net_),
            .in3(N__26355),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.shiftRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(N__36609),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i6_LC_6_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i6_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i6_LC_6_12_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i6_LC_6_12_0  (
            .in0(N__20995),
            .in1(N__22514),
            .in2(_gnd_net_),
            .in3(N__22712),
            .lcout(\Inst_core.Inst_sync.filteredInput_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37543),
            .ce(),
            .sr(N__21080));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3587_1_lut_LC_6_12_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3587_1_lut_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3587_1_lut_LC_6_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3587_1_lut_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20924),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3588_1_lut_LC_6_12_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3588_1_lut_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3588_1_lut_LC_6_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3588_1_lut_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20908),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3589_1_lut_LC_6_12_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3589_1_lut_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3589_1_lut_LC_6_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3589_1_lut_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20897),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3590_1_lut_LC_6_12_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3590_1_lut_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3590_1_lut_LC_6_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3590_1_lut_LC_6_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20980),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3591_1_lut_LC_6_12_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3591_1_lut_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3591_1_lut_LC_6_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3591_1_lut_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20882),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_demux.output_6__12_LC_6_13_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_demux.output_6__12_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_demux.output_6__12_LC_6_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Inst_core.Inst_sync.Inst_demux.output_6__12_LC_6_13_0  (
            .in0(N__23240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.demuxedInput_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i4_LC_6_13_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i4_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i4_LC_6_13_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i4_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__29107),
            .in2(N__31136),
            .in3(N__27360),
            .lcout(divider_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i2_LC_6_13_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i2_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i2_LC_6_13_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i2_LC_6_13_3  (
            .in0(N__31106),
            .in1(N__30909),
            .in2(N__21023),
            .in3(N__31963),
            .lcout(memoryOut_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.i1680_3_lut_4_lut_LC_6_13_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.i1680_3_lut_4_lut_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.i1680_3_lut_4_lut_LC_6_13_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \Inst_core.Inst_sync.i1680_3_lut_4_lut_LC_6_13_4  (
            .in0(N__23239),
            .in1(N__22596),
            .in2(N__21047),
            .in3(N__26380),
            .lcout(),
            .ltout(\Inst_core.Inst_sync.n2789_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i2_LC_6_13_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i2_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i2_LC_6_13_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Inst_core.Inst_sync.output_i2_LC_6_13_5  (
            .in0(N__22920),
            .in1(_gnd_net_),
            .in2(N__21026),
            .in3(N__22804),
            .lcout(syncedInput_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i6_LC_6_13_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i6_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i6_LC_6_13_6 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \Inst_core.Inst_sync.output_i6_LC_6_13_6  (
            .in0(N__22721),
            .in1(N__21010),
            .in2(N__20996),
            .in3(N__22750),
            .lcout(syncedInput_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i4_LC_6_13_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i4_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i4_LC_6_13_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i4_LC_6_13_7  (
            .in0(N__29108),
            .in1(N__22036),
            .in2(_gnd_net_),
            .in3(N__20981),
            .lcout(maskRegister_4_adj_1284),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i5_LC_6_14_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i5_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i5_LC_6_14_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i5_LC_6_14_0  (
            .in0(N__21178),
            .in1(N__22529),
            .in2(_gnd_net_),
            .in3(N__22827),
            .lcout(\Inst_core.Inst_sync.filteredInput_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37569),
            .ce(),
            .sr(N__21059));
    defparam \Inst_core.Inst_sync.Inst_filter.i3478_1_lut_LC_6_14_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3478_1_lut_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3478_1_lut_LC_6_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3478_1_lut_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21109),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4637 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.i3576_1_lut_LC_6_14_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3576_1_lut_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3576_1_lut_LC_6_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3576_1_lut_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20930),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3580_1_lut_LC_6_14_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3580_1_lut_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i3580_1_lut_LC_6_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i3580_1_lut_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20957),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i7_LC_6_15_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i7_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input180Delay_i7_LC_6_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input180Delay_i7_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23111),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input180Delay_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i4_LC_6_15_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i4_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i4_LC_6_15_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i4_LC_6_15_1  (
            .in0(N__31104),
            .in1(N__28027),
            .in2(N__21095),
            .in3(N__31961),
            .lcout(memoryOut_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_demux.output_4__14_LC_6_15_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_demux.output_4__14_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_demux.output_4__14_LC_6_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_demux.output_4__14_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22660),
            .lcout(\Inst_core.Inst_sync.demuxedInput_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7720_LC_6_15_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7720_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7720_LC_6_15_3 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \Inst_core.Inst_sync.n2566_bdd_4_lut_7720_LC_6_15_3  (
            .in0(N__22807),
            .in1(N__22764),
            .in2(N__22832),
            .in3(N__23122),
            .lcout(),
            .ltout(\Inst_core.Inst_sync.n9063_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i5_LC_6_15_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i5_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i5_LC_6_15_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \Inst_core.Inst_sync.output_i5_LC_6_15_4  (
            .in0(N__22766),
            .in1(N__21179),
            .in2(N__21164),
            .in3(N__22894),
            .lcout(syncedInput_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i5_LC_6_15_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i5_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i5_LC_6_15_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i5_LC_6_15_5  (
            .in0(N__31105),
            .in1(N__25455),
            .in2(N__21161),
            .in3(N__31962),
            .lcout(memoryOut_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7679_LC_6_15_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7679_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7679_LC_6_15_6 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \Inst_core.Inst_sync.n2566_bdd_4_lut_7679_LC_6_15_6  (
            .in0(N__22763),
            .in1(N__21144),
            .in2(N__21242),
            .in3(N__22808),
            .lcout(),
            .ltout(\Inst_core.Inst_sync.n9057_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i4_LC_6_15_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i4_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i4_LC_6_15_7 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \Inst_core.Inst_sync.output_i4_LC_6_15_7  (
            .in0(N__21131),
            .in1(N__21110),
            .in2(N__21098),
            .in3(N__22765),
            .lcout(syncedInput_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.i3575_1_lut_LC_6_16_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3575_1_lut_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3575_1_lut_LC_6_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3575_1_lut_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21086),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.i3574_1_lut_LC_6_16_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.i3574_1_lut_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.Inst_filter.i3574_1_lut_LC_6_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.i3574_1_lut_LC_6_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21065),
            .lcout(\Inst_core.Inst_sync.Inst_filter.n4733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i4_LC_6_16_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i4_LC_6_16_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i4_LC_6_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i4_LC_6_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21259),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i4C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.match_84_LC_7_1_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.match_84_LC_7_1_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.match_84_LC_7_1_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.match_84_LC_7_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23642),
            .lcout(\Inst_core.Inst_trigger.stageMatch_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37596),
            .ce(N__32609),
            .sr(N__23411));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i6_LC_7_2_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i6_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i6_LC_7_2_0 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i6_LC_7_2_0  (
            .in0(N__21800),
            .in1(N__21302),
            .in2(N__33557),
            .in3(N__30457),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37585),
            .ce(),
            .sr(N__21227));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i9_4_lut_LC_7_2_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i9_4_lut_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i9_4_lut_LC_7_2_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i9_4_lut_LC_7_2_1  (
            .in0(N__23527),
            .in1(N__23362),
            .in2(N__23573),
            .in3(N__23392),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i15_4_lut_LC_7_2_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i15_4_lut_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i15_4_lut_LC_7_2_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i15_4_lut_LC_7_2_2  (
            .in0(N__21185),
            .in1(N__21206),
            .in2(N__21215),
            .in3(N__21212),
            .lcout(\Inst_core.n31_adj_1174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i11_4_lut_LC_7_2_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i11_4_lut_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i11_4_lut_LC_7_2_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i11_4_lut_LC_7_2_3  (
            .in0(N__23332),
            .in1(N__23821),
            .in2(N__23512),
            .in3(N__23446),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i10_4_lut_LC_7_2_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i10_4_lut_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i10_4_lut_LC_7_2_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i10_4_lut_LC_7_2_4  (
            .in0(N__23803),
            .in1(N__23587),
            .in2(N__23552),
            .in3(N__23491),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i7_LC_7_3_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i7_LC_7_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i7_LC_7_3_0 .LUT_INIT=16'b0011100101101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i7_LC_7_3_0  (
            .in0(N__33538),
            .in1(N__21275),
            .in2(N__21785),
            .in3(N__23053),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37572),
            .ce(),
            .sr(N__21200));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i12_4_lut_LC_7_3_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i12_4_lut_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i12_4_lut_LC_7_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i12_4_lut_LC_7_3_1  (
            .in0(N__23788),
            .in1(N__23473),
            .in2(N__23684),
            .in3(N__23428),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i9_4_lut_LC_7_3_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i9_4_lut_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i9_4_lut_LC_7_3_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i9_4_lut_LC_7_3_2  (
            .in0(N__21448),
            .in1(N__21436),
            .in2(N__21425),
            .in3(N__21400),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i15_4_lut_LC_7_3_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i15_4_lut_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i15_4_lut_LC_7_3_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i15_4_lut_LC_7_3_3  (
            .in0(N__21389),
            .in1(N__21308),
            .in2(N__21377),
            .in3(N__21374),
            .lcout(\Inst_core.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i10_4_lut_LC_7_3_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i10_4_lut_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i10_4_lut_LC_7_3_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i10_4_lut_LC_7_3_4  (
            .in0(N__21358),
            .in1(N__21346),
            .in2(N__21335),
            .in3(N__21319),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i6_LC_7_4_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i6_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i6_LC_7_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i6_LC_7_4_0  (
            .in0(N__36088),
            .in1(N__34424),
            .in2(_gnd_net_),
            .in3(N__21298),
            .lcout(valueRegister_6_adj_1370),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i12_LC_7_4_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i12_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i12_LC_7_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i12_LC_7_4_1  (
            .in0(N__34593),
            .in1(N__29267),
            .in2(_gnd_net_),
            .in3(N__28405),
            .lcout(configRegister_11_adj_1309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i6_LC_7_4_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i6_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i6_LC_7_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i6_LC_7_4_2  (
            .in0(N__31402),
            .in1(N__21286),
            .in2(_gnd_net_),
            .in3(N__26088),
            .lcout(configRegister_5_adj_1395),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i11_LC_7_4_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i11_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i11_LC_7_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i11_LC_7_4_3  (
            .in0(N__35799),
            .in1(N__25588),
            .in2(_gnd_net_),
            .in3(N__23458),
            .lcout(configRegister_10_adj_1350),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i11_LC_7_4_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i11_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i11_LC_7_4_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i11_LC_7_4_4  (
            .in0(N__25587),
            .in1(N__34594),
            .in2(N__34840),
            .in3(N__35068),
            .lcout(cmd_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i7_LC_7_4_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i7_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i7_LC_7_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i7_LC_7_4_5  (
            .in0(N__36089),
            .in1(N__27198),
            .in2(_gnd_net_),
            .in3(N__21274),
            .lcout(valueRegister_7_adj_1369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i12_LC_7_4_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i12_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i12_LC_7_4_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i12_LC_7_4_6  (
            .in0(N__34595),
            .in1(N__26087),
            .in2(_gnd_net_),
            .in3(N__21517),
            .lcout(configRegister_11_adj_1389),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i11_LC_7_4_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i11_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i11_LC_7_4_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i11_LC_7_4_7  (
            .in0(N__26086),
            .in1(N__25589),
            .in2(_gnd_net_),
            .in3(N__21505),
            .lcout(configRegister_10_adj_1390),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i0_LC_7_5_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i0_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i0_LC_7_5_0 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i0_LC_7_5_0  (
            .in0(N__26342),
            .in1(N__21473),
            .in2(N__21494),
            .in3(N__21755),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i1_LC_7_5_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i1_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i1_LC_7_5_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i1_LC_7_5_1  (
            .in0(N__21472),
            .in1(N__31701),
            .in2(_gnd_net_),
            .in3(N__26335),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i2_LC_7_5_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i2_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i2_LC_7_5_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i2_LC_7_5_2  (
            .in0(N__26336),
            .in1(N__33456),
            .in2(N__31708),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i3_LC_7_5_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i3_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i3_LC_7_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i3_LC_7_5_3  (
            .in0(N__33457),
            .in1(N__28635),
            .in2(_gnd_net_),
            .in3(N__26337),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i4_LC_7_5_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i4_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i4_LC_7_5_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i4_LC_7_5_4  (
            .in0(N__26338),
            .in1(_gnd_net_),
            .in2(N__28642),
            .in3(N__32373),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i5_LC_7_5_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i5_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i5_LC_7_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i5_LC_7_5_5  (
            .in0(N__32374),
            .in1(N__28113),
            .in2(_gnd_net_),
            .in3(N__26339),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i6_LC_7_5_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i6_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i6_LC_7_5_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i6_LC_7_5_6  (
            .in0(N__26340),
            .in1(_gnd_net_),
            .in2(N__28120),
            .in3(N__25527),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i7_LC_7_5_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i7_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i7_LC_7_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_i0_i7_LC_7_5_7  (
            .in0(N__25528),
            .in1(N__21796),
            .in2(_gnd_net_),
            .in3(N__26341),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.shiftRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(N__36643),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i4_LC_7_6_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i4_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i4_LC_7_6_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i4_LC_7_6_0  (
            .in0(N__35060),
            .in1(N__26652),
            .in2(N__29128),
            .in3(N__34796),
            .lcout(cmd_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i16_LC_7_6_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i16_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i16_LC_7_6_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i16_LC_7_6_1  (
            .in0(N__33913),
            .in1(N__26076),
            .in2(_gnd_net_),
            .in3(N__21766),
            .lcout(configRegister_15_adj_1385),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i9_LC_7_6_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i9_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i9_LC_7_6_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i9_LC_7_6_3  (
            .in0(N__23978),
            .in1(_gnd_net_),
            .in2(N__28489),
            .in3(N__29333),
            .lcout(configRegister_8_adj_1312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i23_LC_7_6_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i23_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i23_LC_7_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i23_LC_7_6_4  (
            .in0(N__26075),
            .in1(N__21754),
            .in2(_gnd_net_),
            .in3(N__22219),
            .lcout(configRegister_24_adj_1378),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i5_LC_7_6_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i5_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i5_LC_7_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i5_LC_7_6_5  (
            .in0(N__23917),
            .in1(N__31352),
            .in2(_gnd_net_),
            .in3(N__25639),
            .lcout(maskRegister_5_adj_1363),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.disabledGroupsReg_i0_i0_LC_7_6_6 .C_ON=1'b0;
    defparam \Inst_eia232.disabledGroupsReg_i0_i0_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.disabledGroupsReg_i0_i0_LC_7_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_eia232.disabledGroupsReg_i0_i0_LC_7_6_6  (
            .in0(N__22285),
            .in1(N__29676),
            .in2(_gnd_net_),
            .in3(N__21547),
            .lcout(disabledGroupsReg_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i0_LC_7_6_7 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i0_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_transmitter.disabledBuffer_i0_LC_7_6_7 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \Inst_eia232.Inst_transmitter.disabledBuffer_i0_LC_7_6_7  (
            .in0(N__21731),
            .in1(N__21681),
            .in2(N__21551),
            .in3(N__21532),
            .lcout(\Inst_eia232.Inst_transmitter.disabledBuffer_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i24_LC_7_7_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i24_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i24_LC_7_7_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i24_LC_7_7_0  (
            .in0(N__35050),
            .in1(N__22203),
            .in2(N__29756),
            .in3(N__34801),
            .lcout(cmd_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i1_LC_7_7_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i1_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i1_LC_7_7_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i1_LC_7_7_1  (
            .in0(N__34206),
            .in1(N__34800),
            .in2(N__35954),
            .in3(N__35051),
            .lcout(cmd_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i14_LC_7_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i14_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i14_LC_7_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i14_LC_7_7_2  (
            .in0(N__29383),
            .in1(N__34106),
            .in2(_gnd_net_),
            .in3(N__33835),
            .lcout(configRegister_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i6_LC_7_7_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i6_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i6_LC_7_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i6_LC_7_7_3  (
            .in0(N__29457),
            .in1(N__34410),
            .in2(_gnd_net_),
            .in3(N__27394),
            .lcout(valueRegister_6_adj_1330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i14_LC_7_7_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i14_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i14_LC_7_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i14_LC_7_7_4  (
            .in0(N__29384),
            .in1(N__29332),
            .in2(_gnd_net_),
            .in3(N__28804),
            .lcout(configRegister_13_adj_1307),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i21_LC_7_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i21_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i21_LC_7_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i21_LC_7_7_5  (
            .in0(N__24175),
            .in1(N__26102),
            .in2(_gnd_net_),
            .in3(N__21925),
            .lcout(configRegister_22_adj_1380),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i22_LC_7_7_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i22_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i22_LC_7_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i22_LC_7_7_6  (
            .in0(N__29745),
            .in1(N__34107),
            .in2(_gnd_net_),
            .in3(N__21904),
            .lcout(configRegister_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i8_LC_7_7_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i8_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i8_LC_7_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i8_LC_7_7_7  (
            .in0(N__31197),
            .in1(N__23985),
            .in2(_gnd_net_),
            .in3(N__27262),
            .lcout(divider_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i8_LC_7_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i8_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i8_LC_7_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i8_LC_7_8_0  (
            .in0(N__35476),
            .in1(N__23997),
            .in2(_gnd_net_),
            .in3(N__24265),
            .lcout(bwd_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i0_LC_7_8_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i0_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i0_LC_7_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.maskRegister_i0_i0_LC_7_8_1  (
            .in0(N__21890),
            .in1(N__35925),
            .in2(_gnd_net_),
            .in3(N__21830),
            .lcout(maskRegister_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i19_LC_7_8_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i19_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i19_LC_7_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i19_LC_7_8_2  (
            .in0(N__26112),
            .in1(N__26536),
            .in2(_gnd_net_),
            .in3(N__21816),
            .lcout(configRegister_20_adj_1382),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i21_LC_7_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i21_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i21_LC_7_8_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i21_LC_7_8_3  (
            .in0(N__24153),
            .in1(N__35795),
            .in2(_gnd_net_),
            .in3(N__22102),
            .lcout(configRegister_22_adj_1340),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i25_LC_7_8_5 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i25_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i25_LC_7_8_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i25_LC_7_8_5  (
            .in0(N__34797),
            .in1(N__24101),
            .in2(N__22216),
            .in3(N__34959),
            .lcout(cmd_32),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i30_LC_7_8_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i30_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i30_LC_7_8_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i30_LC_7_8_6  (
            .in0(N__34958),
            .in1(N__24061),
            .in2(N__24390),
            .in3(N__34798),
            .lcout(cmd_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i11_LC_7_8_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i11_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i11_LC_7_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i11_LC_7_8_7  (
            .in0(N__34582),
            .in1(N__31196),
            .in2(_gnd_net_),
            .in3(N__30771),
            .lcout(divider_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i20_LC_7_9_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i20_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i20_LC_7_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i20_LC_7_9_0  (
            .in0(N__22061),
            .in1(N__24668),
            .in2(_gnd_net_),
            .in3(N__34084),
            .lcout(configRegister_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i6_LC_7_9_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i6_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i6_LC_7_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.maskRegister_i0_i6_LC_7_9_1  (
            .in0(N__22024),
            .in1(N__34422),
            .in2(_gnd_net_),
            .in3(N__29779),
            .lcout(maskRegister_6_adj_1282),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i1_LC_7_9_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i1_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i1_LC_7_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i1_LC_7_9_2  (
            .in0(N__34527),
            .in1(N__34231),
            .in2(_gnd_net_),
            .in3(N__22135),
            .lcout(valueRegister_1_adj_1295),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i9_LC_7_9_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i9_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i9_LC_7_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i9_LC_7_9_3  (
            .in0(N__26586),
            .in1(N__31185),
            .in2(_gnd_net_),
            .in3(N__24888),
            .lcout(divider_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i20_LC_7_9_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i20_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i20_LC_7_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i20_LC_7_9_4  (
            .in0(N__35820),
            .in1(N__24669),
            .in2(_gnd_net_),
            .in3(N__21952),
            .lcout(configRegister_21_adj_1341),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i16_LC_7_9_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i16_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i16_LC_7_9_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i16_LC_7_9_6  (
            .in0(N__35017),
            .in1(N__33898),
            .in2(N__36184),
            .in3(N__34804),
            .lcout(cmd_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_flags.inverted_18_LC_7_9_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_flags.inverted_18_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_flags.inverted_18_LC_7_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_flags.inverted_18_LC_7_9_7  (
            .in0(N__22615),
            .in1(N__27191),
            .in2(_gnd_net_),
            .in3(N__22278),
            .lcout(flagInverted),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i8_LC_7_10_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i8_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i8_LC_7_10_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i8_LC_7_10_0  (
            .in0(N__22217),
            .in1(N__35406),
            .in2(_gnd_net_),
            .in3(N__24436),
            .lcout(fwd_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i11_LC_7_10_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i11_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i11_LC_7_10_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i11_LC_7_10_1  (
            .in0(N__28177),
            .in1(_gnd_net_),
            .in2(N__35441),
            .in3(N__24251),
            .lcout(fwd_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i5_LC_7_10_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i5_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i5_LC_7_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i5_LC_7_10_2  (
            .in0(N__35407),
            .in1(N__24685),
            .in2(_gnd_net_),
            .in3(N__22346),
            .lcout(fwd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i20_LC_7_10_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i20_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i20_LC_7_10_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i20_LC_7_10_3  (
            .in0(N__31164),
            .in1(_gnd_net_),
            .in2(N__26534),
            .in3(N__25050),
            .lcout(divider_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i5_LC_7_10_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i5_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i5_LC_7_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i5_LC_7_10_4  (
            .in0(N__31351),
            .in1(N__35401),
            .in2(_gnd_net_),
            .in3(N__26785),
            .lcout(bwd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i6_LC_7_10_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i6_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i6_LC_7_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i6_LC_7_10_5  (
            .in0(N__35405),
            .in1(N__24176),
            .in2(_gnd_net_),
            .in3(N__22361),
            .lcout(fwd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i22_LC_7_10_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i22_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i22_LC_7_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i22_LC_7_10_6  (
            .in0(N__24177),
            .in1(N__31165),
            .in2(_gnd_net_),
            .in3(N__32046),
            .lcout(divider_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i19_LC_7_10_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i19_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i19_LC_7_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i19_LC_7_10_7  (
            .in0(N__26524),
            .in1(N__34120),
            .in2(_gnd_net_),
            .in3(N__22161),
            .lcout(configRegister_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i1_LC_7_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i1_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i1_LC_7_11_0 .LUT_INIT=16'b0110011001011010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i1_LC_7_11_0  (
            .in0(N__22142),
            .in1(N__22124),
            .in2(N__33645),
            .in3(N__30359),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37545),
            .ce(),
            .sr(N__22400));
    defparam \Inst_core.Inst_controller.i10_4_lut_LC_7_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i10_4_lut_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i10_4_lut_LC_7_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_controller.i10_4_lut_LC_7_11_1  (
            .in0(N__24449),
            .in1(N__24185),
            .in2(N__30173),
            .in3(N__24470),
            .lcout(),
            .ltout(\Inst_core.Inst_controller.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_55_LC_7_11_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_55_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_55_LC_7_11_2 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \Inst_core.Inst_controller.i1_4_lut_adj_55_LC_7_11_2  (
            .in0(N__37663),
            .in1(N__22382),
            .in2(N__22364),
            .in3(N__24218),
            .lcout(),
            .ltout(\Inst_core.Inst_controller.n4_adj_986_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_56_LC_7_11_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_56_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_56_LC_7_11_3 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \Inst_core.Inst_controller.i1_4_lut_adj_56_LC_7_11_3  (
            .in0(N__22360),
            .in1(N__36989),
            .in2(N__22349),
            .in3(N__22331),
            .lcout(),
            .ltout(\Inst_core.Inst_controller.n4_adj_987_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_57_LC_7_11_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_57_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_57_LC_7_11_4 .LUT_INIT=16'b1111011011111111;
    LogicCell40 \Inst_core.Inst_controller.i1_4_lut_adj_57_LC_7_11_4  (
            .in0(N__37025),
            .in1(N__22345),
            .in2(N__22334),
            .in3(N__29861),
            .lcout(\Inst_core.Inst_controller.nstate_1_N_829_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i15_2_lut_LC_7_11_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i15_2_lut_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i15_2_lut_LC_7_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Inst_core.Inst_controller.i15_2_lut_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__24035),
            .in2(_gnd_net_),
            .in3(N__37697),
            .lcout(\Inst_core.Inst_controller.n8486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i3_LC_7_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i3_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i3_LC_7_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_sync.output_i3_LC_7_12_0  (
            .in0(N__22801),
            .in1(N__22849),
            .in2(_gnd_net_),
            .in3(N__22421),
            .lcout(syncedInput_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i0_LC_7_12_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i0_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i0_LC_7_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_sync.output_i0_LC_7_12_1  (
            .in0(N__22325),
            .in1(N__22802),
            .in2(_gnd_net_),
            .in3(N__22622),
            .lcout(syncedInput_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i5_LC_7_12_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i5_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i5_LC_7_12_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i5_LC_7_12_2  (
            .in0(N__29482),
            .in1(N__24823),
            .in2(_gnd_net_),
            .in3(N__31370),
            .lcout(valueRegister_5_adj_1331),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i7_LC_7_12_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i7_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i7_LC_7_12_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i7_LC_7_12_3  (
            .in0(N__22477),
            .in1(N__29483),
            .in2(_gnd_net_),
            .in3(N__27199),
            .lcout(valueRegister_7_adj_1329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i0_LC_7_12_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i0_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i0_LC_7_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i0_LC_7_12_5  (
            .in0(N__27050),
            .in1(N__35984),
            .in2(_gnd_net_),
            .in3(N__26902),
            .lcout(maskRegister_0_adj_1328),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i3_LC_7_12_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i3_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i3_LC_7_12_6 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i3_LC_7_12_6  (
            .in0(N__31163),
            .in1(N__32313),
            .in2(N__22502),
            .in3(N__31955),
            .lcout(memoryOut_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i7_LC_7_12_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i7_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i7_LC_7_12_7 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \Inst_core.Inst_sync.output_i7_LC_7_12_7  (
            .in0(N__22951),
            .in1(N__22751),
            .in2(N__26969),
            .in3(N__22874),
            .lcout(syncedInput_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i7_LC_7_13_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i7_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i7_LC_7_13_0 .LUT_INIT=16'b0011100101101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i7_LC_7_13_0  (
            .in0(N__35612),
            .in1(N__22478),
            .in2(N__25106),
            .in3(N__23036),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37571),
            .ce(),
            .sr(N__26456));
    defparam \Inst_core.Inst_sampler.i7222_4_lut_LC_7_13_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7222_4_lut_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7222_4_lut_LC_7_13_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_sampler.i7222_4_lut_LC_7_13_1  (
            .in0(N__25054),
            .in1(N__27854),
            .in2(N__32056),
            .in3(N__27806),
            .lcout(\Inst_core.Inst_sampler.n8590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7234_4_lut_LC_7_13_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7234_4_lut_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7234_4_lut_LC_7_13_2 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_sampler.i7234_4_lut_LC_7_13_2  (
            .in0(N__31655),
            .in1(N__24871),
            .in2(N__24899),
            .in3(N__27506),
            .lcout(\Inst_core.Inst_sampler.n8602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.i1678_3_lut_4_lut_LC_7_13_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.i1678_3_lut_4_lut_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.i1678_3_lut_4_lut_LC_7_13_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \Inst_core.Inst_sync.i1678_3_lut_4_lut_LC_7_13_3  (
            .in0(N__22600),
            .in1(N__26359),
            .in2(N__22466),
            .in3(N__23276),
            .lcout(\Inst_core.Inst_sync.n2787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.i5524_1_lut_2_lut_LC_7_13_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.i5524_1_lut_2_lut_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.i5524_1_lut_2_lut_LC_7_13_4 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \Inst_core.Inst_sync.i5524_1_lut_2_lut_LC_7_13_4  (
            .in0(N__26358),
            .in1(N__22599),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.n2564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.i1682_3_lut_4_lut_LC_7_13_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.i1682_3_lut_4_lut_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.i1682_3_lut_4_lut_LC_7_13_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \Inst_core.Inst_sync.i1682_3_lut_4_lut_LC_7_13_5  (
            .in0(N__23204),
            .in1(N__22598),
            .in2(N__22442),
            .in3(N__26360),
            .lcout(\Inst_core.Inst_sync.n2791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.i1684_3_lut_4_lut_LC_7_13_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.i1684_3_lut_4_lut_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.i1684_3_lut_4_lut_LC_7_13_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \Inst_core.Inst_sync.i1684_3_lut_4_lut_LC_7_13_6  (
            .in0(N__26361),
            .in1(N__22601),
            .in2(N__22646),
            .in3(N__22661),
            .lcout(\Inst_core.Inst_sync.n2793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.i1459_3_lut_LC_7_13_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.i1459_3_lut_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.i1459_3_lut_LC_7_13_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \Inst_core.Inst_sync.i1459_3_lut_LC_7_13_7  (
            .in0(N__22616),
            .in1(N__22597),
            .in2(_gnd_net_),
            .in3(N__26357),
            .lcout(\Inst_core.Inst_sync.n2566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.output_i1_LC_7_14_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.output_i1_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.output_i1_LC_7_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_sync.output_i1_LC_7_14_0  (
            .in0(N__22559),
            .in1(N__22803),
            .in2(_gnd_net_),
            .in3(N__22535),
            .lcout(syncedInput_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i5_LC_7_14_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i5_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i5_LC_7_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i5_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22828),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i6_LC_7_14_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i6_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i6_LC_7_14_2 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i6_LC_7_14_2  (
            .in0(N__31138),
            .in1(N__30405),
            .in2(N__22523),
            .in3(N__31949),
            .lcout(memoryOut_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i15_LC_7_14_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i15_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i15_LC_7_14_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i15_LC_7_14_3  (
            .in0(N__33914),
            .in1(N__31140),
            .in2(_gnd_net_),
            .in3(N__24803),
            .lcout(divider_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i6_LC_7_14_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i6_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i6_LC_7_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i6_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22711),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i16_LC_7_14_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i16_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i16_LC_7_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i16_LC_7_14_6  (
            .in0(N__31137),
            .in1(N__36185),
            .in2(_gnd_net_),
            .in3(N__24749),
            .lcout(divider_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i0_LC_7_14_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i0_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i0_LC_7_14_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i0_LC_7_14_7  (
            .in0(N__35997),
            .in1(N__31139),
            .in2(_gnd_net_),
            .in3(N__31567),
            .lcout(divider_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_demux.output_7__11_LC_7_15_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_demux.output_7__11_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_demux.output_7__11_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_demux.output_7__11_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23203),
            .lcout(\Inst_core.Inst_sync.demuxedInput_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i2_LC_7_15_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i2_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i2_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i2_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23261),
            .lcout(\Inst_core.Inst_sync.demuxedInput_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_demux.output_5__13_LC_7_15_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_demux.output_5__13_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_demux.output_5__13_LC_7_15_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Inst_core.Inst_sync.Inst_demux.output_5__13_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__23275),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.demuxedInput_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7729_LC_7_15_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7729_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_7729_LC_7_15_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \Inst_core.Inst_sync.n2566_bdd_4_lut_7729_LC_7_15_3  (
            .in0(N__22752),
            .in1(N__22806),
            .in2(N__31435),
            .in3(N__23110),
            .lcout(\Inst_core.Inst_sync.n9117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i3_LC_7_15_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i3_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i3_LC_7_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i3_LC_7_15_4  (
            .in0(N__23228),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.demuxedInput_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i5_LC_7_15_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i5_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i5_LC_7_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i5_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23150),
            .lcout(\Inst_core.Inst_sync.synchronizedInput_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_LC_7_15_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sync.n2566_bdd_4_lut_LC_7_15_6 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \Inst_core.Inst_sync.n2566_bdd_4_lut_LC_7_15_6  (
            .in0(N__22805),
            .in1(N__22753),
            .in2(N__22707),
            .in3(N__23161),
            .lcout(\Inst_core.Inst_sync.n9129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i6_LC_7_15_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i6_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i6_LC_7_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i6_LC_7_15_7  (
            .in0(N__23189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.synchronizedInput_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i0_LC_7_16_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i0_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i0_LC_7_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i0_LC_7_16_0  (
            .in0(N__22681),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i1_LC_7_16_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i1_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i1_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i1_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23303),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i2_LC_7_16_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i2_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i2_LC_7_16_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i2_LC_7_16_2  (
            .in0(N__23257),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i3_LC_7_16_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i3_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i3_LC_7_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i3_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23227),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i6_LC_7_16_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i6_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i6_LC_7_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i6_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23188),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i5_LC_7_16_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i5_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i5_LC_7_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i5_LC_7_16_5  (
            .in0(N__23149),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput180_i7_LC_7_16_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i7_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput180_i7_LC_7_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput180_i7_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31459),
            .lcout(\Inst_core.Inst_sync.synchronizedInput180_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVInst_core.Inst_sync.synchronizedInput180_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_2_lut_LC_8_1_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_2_lut_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_2_lut_LC_8_1_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_2_lut_LC_8_1_0  (
            .in0(N__36635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25226),
            .lcout(\Inst_core.n8518 ),
            .ltout(\Inst_core.n8518_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_decoder.i17_4_lut_LC_8_1_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.i17_4_lut_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_decoder.i17_4_lut_LC_8_1_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Inst_core.Inst_decoder.i17_4_lut_LC_8_1_1  (
            .in0(N__23641),
            .in1(N__32503),
            .in2(N__23099),
            .in3(N__32602),
            .lcout(\Inst_core.Inst_decoder.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i7_LC_8_1_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i7_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i7_LC_8_1_2 .LUT_INIT=16'b0101100101101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i7_LC_8_1_2  (
            .in0(N__23096),
            .in1(N__30345),
            .in2(N__23078),
            .in3(N__23054),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37607),
            .ce(),
            .sr(N__26918));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i7501_2_lut_LC_8_1_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i7501_2_lut_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i7501_2_lut_LC_8_1_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i7501_2_lut_LC_8_1_3  (
            .in0(N__25227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36634),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n8808_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_4_lut_adj_73_LC_8_1_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_4_lut_adj_73_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_4_lut_adj_73_LC_8_1_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i1_4_lut_adj_73_LC_8_1_4  (
            .in0(N__25241),
            .in1(N__36854),
            .in2(N__23414),
            .in3(N__25183),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i7621_2_lut_3_lut_4_lut_LC_8_1_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i7621_2_lut_3_lut_4_lut_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i7621_2_lut_3_lut_4_lut_LC_8_1_5 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i7621_2_lut_3_lut_4_lut_LC_8_1_5  (
            .in0(N__25228),
            .in1(N__36636),
            .in2(N__36873),
            .in3(N__25184),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i2_3_lut_LC_8_1_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i2_3_lut_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i2_3_lut_LC_8_1_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Inst_core.Inst_sampler.i2_3_lut_LC_8_1_6  (
            .in0(N__36633),
            .in1(N__25182),
            .in2(_gnd_net_),
            .in3(N__25225),
            .lcout(\Inst_core.n1639 ),
            .ltout(\Inst_core.n1639_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7669_1_lut_LC_8_1_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7669_1_lut_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7669_1_lut_LC_8_1_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \Inst_core.Inst_sampler.i7669_1_lut_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23405),
            .in3(_gnd_net_),
            .lcout(\Inst_core.n9054 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i0_LC_8_2_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i0_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i0_LC_8_2_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i0_LC_8_2_0  (
            .in0(N__28136),
            .in1(N__23402),
            .in2(N__23396),
            .in3(N__23381),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_0 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7899 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i1_LC_8_2_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i1_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i1_LC_8_2_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i1_LC_8_2_1  (
            .in0(N__23378),
            .in1(N__23363),
            .in2(N__23770),
            .in3(N__23351),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_1 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7899 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7900 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i2_LC_8_2_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i2_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i2_LC_8_2_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i2_LC_8_2_2  (
            .in0(N__23348),
            .in1(N__23333),
            .in2(N__23751),
            .in3(N__23321),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_2 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7900 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7901 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i3_LC_8_2_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i3_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i3_LC_8_2_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i3_LC_8_2_3  (
            .in0(N__23318),
            .in1(N__23721),
            .in2(N__23591),
            .in3(N__23576),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_3 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7901 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7902 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i4_LC_8_2_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i4_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i4_LC_8_2_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i4_LC_8_2_4  (
            .in0(N__25658),
            .in1(N__23569),
            .in2(N__23752),
            .in3(N__23555),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_4 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7902 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7903 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i5_LC_8_2_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i5_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i5_LC_8_2_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i5_LC_8_2_5  (
            .in0(N__23867),
            .in1(N__23725),
            .in2(N__23551),
            .in3(N__23531),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_5 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7903 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7904 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i6_LC_8_2_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i6_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i6_LC_8_2_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i6_LC_8_2_6  (
            .in0(N__24353),
            .in1(N__23528),
            .in2(N__23753),
            .in3(N__23516),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_6 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7904 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7905 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i7_LC_8_2_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i7_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i7_LC_8_2_7 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i7_LC_8_2_7  (
            .in0(N__23618),
            .in1(N__23729),
            .in2(N__23513),
            .in3(N__23495),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_7 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7905 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7906 ),
            .clk(N__37598),
            .ce(N__23669),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i8_LC_8_3_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i8_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i8_LC_8_3_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i8_LC_8_3_0  (
            .in0(N__24017),
            .in1(N__23492),
            .in2(N__23771),
            .in3(N__23480),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_8 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7907 ),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i9_LC_8_3_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i9_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i9_LC_8_3_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i9_LC_8_3_1  (
            .in0(N__23837),
            .in1(N__23757),
            .in2(N__23477),
            .in3(N__23462),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_9 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7907 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7908 ),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i10_LC_8_3_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i10_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i10_LC_8_3_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i10_LC_8_3_2  (
            .in0(N__23459),
            .in1(N__23447),
            .in2(N__23772),
            .in3(N__23435),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_10 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7908 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7909 ),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i11_LC_8_3_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i11_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i11_LC_8_3_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i11_LC_8_3_3  (
            .in0(N__23603),
            .in1(N__23761),
            .in2(N__23432),
            .in3(N__23417),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_11 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7909 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7910 ),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i12_LC_8_3_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i12_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i12_LC_8_3_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i12_LC_8_3_4  (
            .in0(N__25955),
            .in1(N__23822),
            .in2(N__23773),
            .in3(N__23810),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_12 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7910 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7911 ),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i13_LC_8_3_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i13_LC_8_3_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i13_LC_8_3_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i13_LC_8_3_5  (
            .in0(N__25562),
            .in1(N__23765),
            .in2(N__23807),
            .in3(N__23792),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_13 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7911 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7912 ),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i14_LC_8_3_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i14_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i14_LC_8_3_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i14_LC_8_3_6  (
            .in0(N__23852),
            .in1(N__23789),
            .in2(N__23774),
            .in3(N__23777),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_14 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7912 ),
            .carryout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7913 ),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i15_LC_8_3_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i15_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i15_LC_8_3_7 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.counter__i15_LC_8_3_7  (
            .in0(N__23769),
            .in1(N__23683),
            .in2(N__23939),
            .in3(N__23687),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37587),
            .ce(N__23668),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i25_LC_8_4_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i25_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i25_LC_8_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i25_LC_8_4_0  (
            .in0(N__23640),
            .in1(N__28178),
            .in2(_gnd_net_),
            .in3(N__35856),
            .lcout(\Inst_core.configRegister_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i14_LC_8_4_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i14_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i14_LC_8_4_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i14_LC_8_4_1  (
            .in0(N__29354),
            .in1(N__34810),
            .in2(N__30119),
            .in3(N__35069),
            .lcout(cmd_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i8_LC_8_4_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i8_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i8_LC_8_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i8_LC_8_4_2  (
            .in0(N__27197),
            .in1(N__23614),
            .in2(_gnd_net_),
            .in3(N__35857),
            .lcout(configRegister_7_adj_1353),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i12_LC_8_4_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i12_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i12_LC_8_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i12_LC_8_4_3  (
            .in0(N__35854),
            .in1(N__34591),
            .in2(_gnd_net_),
            .in3(N__23602),
            .lcout(configRegister_11_adj_1349),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i13_LC_8_4_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i13_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i13_LC_8_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i13_LC_8_4_4  (
            .in0(N__26136),
            .in1(N__35308),
            .in2(_gnd_net_),
            .in3(N__23878),
            .lcout(configRegister_12_adj_1388),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i6_LC_8_4_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i6_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i6_LC_8_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i6_LC_8_4_5  (
            .in0(N__35855),
            .in1(N__31374),
            .in2(_gnd_net_),
            .in3(N__23863),
            .lcout(configRegister_5_adj_1355),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i3_LC_8_4_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i3_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i3_LC_8_4_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i3_LC_8_4_6  (
            .in0(N__32749),
            .in1(N__34121),
            .in2(_gnd_net_),
            .in3(N__29678),
            .lcout(configRegister_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i3_LC_8_4_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i3_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i3_LC_8_4_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i3_LC_8_4_7  (
            .in0(N__36104),
            .in1(N__26698),
            .in2(_gnd_net_),
            .in3(N__32392),
            .lcout(valueRegister_3_adj_1373),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i4_LC_8_5_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i4_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i4_LC_8_5_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i4_LC_8_5_0  (
            .in0(N__34123),
            .in1(N__32719),
            .in2(_gnd_net_),
            .in3(N__26654),
            .lcout(configRegister_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i15_LC_8_5_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i15_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i15_LC_8_5_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i15_LC_8_5_1  (
            .in0(N__35852),
            .in1(N__30114),
            .in2(_gnd_net_),
            .in3(N__23848),
            .lcout(configRegister_14_adj_1346),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i11_LC_8_5_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i11_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i11_LC_8_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i11_LC_8_5_2  (
            .in0(N__34122),
            .in1(N__25593),
            .in2(_gnd_net_),
            .in3(N__33076),
            .lcout(configRegister_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i13_LC_8_5_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i13_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i13_LC_8_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i13_LC_8_5_3  (
            .in0(N__29310),
            .in1(N__35307),
            .in2(_gnd_net_),
            .in3(N__28372),
            .lcout(configRegister_12_adj_1308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i10_LC_8_5_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i10_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i10_LC_8_5_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i10_LC_8_5_5  (
            .in0(N__23833),
            .in1(N__35813),
            .in2(_gnd_net_),
            .in3(N__26597),
            .lcout(configRegister_9_adj_1351),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i8_LC_8_5_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i8_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i8_LC_8_5_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i8_LC_8_5_6  (
            .in0(N__29311),
            .in1(N__28507),
            .in2(_gnd_net_),
            .in3(N__27192),
            .lcout(configRegister_7_adj_1313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i9_LC_8_5_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i9_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i9_LC_8_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i9_LC_8_5_7  (
            .in0(N__35853),
            .in1(N__24010),
            .in2(_gnd_net_),
            .in3(N__23999),
            .lcout(configRegister_8_adj_1352),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i18_LC_8_6_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i18_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i18_LC_8_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i18_LC_8_6_0  (
            .in0(N__29555),
            .in1(N__35851),
            .in2(_gnd_net_),
            .in3(N__28927),
            .lcout(configRegister_17_adj_1343),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i9_LC_8_6_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i9_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i9_LC_8_6_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i9_LC_8_6_1  (
            .in0(N__34095),
            .in1(N__33130),
            .in2(_gnd_net_),
            .in3(N__23993),
            .lcout(configRegister_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i8_LC_8_6_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i8_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i8_LC_8_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i8_LC_8_6_2  (
            .in0(N__34085),
            .in1(N__33163),
            .in2(_gnd_net_),
            .in3(N__27174),
            .lcout(configRegister_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i1_LC_8_6_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i1_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i1_LC_8_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i1_LC_8_6_3  (
            .in0(N__23919),
            .in1(N__34237),
            .in2(_gnd_net_),
            .in3(N__26426),
            .lcout(maskRegister_1_adj_1367),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i17_LC_8_6_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i17_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i17_LC_8_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i17_LC_8_6_4  (
            .in0(N__29554),
            .in1(N__31198),
            .in2(_gnd_net_),
            .in3(N__27237),
            .lcout(divider_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i16_LC_8_6_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i16_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i16_LC_8_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i16_LC_8_6_5  (
            .in0(N__35850),
            .in1(N__33928),
            .in2(_gnd_net_),
            .in3(N__23932),
            .lcout(configRegister_15_adj_1345),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i0_LC_8_6_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i0_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i0_LC_8_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i0_LC_8_6_6  (
            .in0(N__26441),
            .in1(N__35928),
            .in2(_gnd_net_),
            .in3(N__23918),
            .lcout(maskRegister_0_adj_1368),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i2_LC_8_6_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i2_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i2_LC_8_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.maskRegister_i0_i2_LC_8_6_7  (
            .in0(N__23920),
            .in1(N__29677),
            .in2(_gnd_net_),
            .in3(N__26414),
            .lcout(maskRegister_2_adj_1366),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i11_LC_8_7_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i11_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i11_LC_8_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i11_LC_8_7_0  (
            .in0(N__29330),
            .in1(N__25609),
            .in2(_gnd_net_),
            .in3(N__28426),
            .lcout(configRegister_10_adj_1310),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i6_LC_8_7_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i6_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i6_LC_8_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i6_LC_8_7_1  (
            .in0(N__27053),
            .in1(N__34420),
            .in2(_gnd_net_),
            .in3(N__25868),
            .lcout(maskRegister_6_adj_1322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i13_LC_8_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i13_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i13_LC_8_7_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i13_LC_8_7_2  (
            .in0(N__29382),
            .in1(_gnd_net_),
            .in2(N__31199),
            .in3(N__24771),
            .lcout(divider_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i5_LC_8_7_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i5_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i5_LC_8_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i5_LC_8_7_3  (
            .in0(N__27052),
            .in1(N__31364),
            .in2(_gnd_net_),
            .in3(N__25895),
            .lcout(maskRegister_5_adj_1323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i10_LC_8_7_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i10_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i10_LC_8_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i10_LC_8_7_4  (
            .in0(N__26585),
            .in1(N__26120),
            .in2(_gnd_net_),
            .in3(N__24073),
            .lcout(configRegister_9_adj_1391),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i24_LC_8_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i24_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i24_LC_8_7_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i24_LC_8_7_5  (
            .in0(N__35671),
            .in1(_gnd_net_),
            .in2(N__26135),
            .in3(N__33514),
            .lcout(configRegister_26_adj_1377),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i10_LC_8_7_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i10_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i10_LC_8_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i10_LC_8_7_6  (
            .in0(N__35444),
            .in1(N__25608),
            .in2(_gnd_net_),
            .in3(N__24463),
            .lcout(bwd_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i14_LC_8_7_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i14_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i14_LC_8_7_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i14_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__31192),
            .in2(N__30113),
            .in3(N__24711),
            .lcout(divider_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i14_LC_8_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i14_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i14_LC_8_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i14_LC_8_8_0  (
            .in0(N__24062),
            .in1(N__24034),
            .in2(_gnd_net_),
            .in3(N__35478),
            .lcout(\Inst_core.Inst_controller.fwd_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i23_LC_8_8_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i23_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i23_LC_8_8_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i23_LC_8_8_1  (
            .in0(N__34960),
            .in1(N__29752),
            .in2(N__24168),
            .in3(N__34789),
            .lcout(cmd_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i10_LC_8_8_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i10_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i10_LC_8_8_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i10_LC_8_8_2  (
            .in0(N__26584),
            .in1(N__34961),
            .in2(N__25613),
            .in3(N__34802),
            .lcout(cmd_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i18_LC_8_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i18_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i18_LC_8_8_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i18_LC_8_8_3  (
            .in0(N__29541),
            .in1(N__26127),
            .in2(_gnd_net_),
            .in3(N__25801),
            .lcout(configRegister_17_adj_1383),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i26_LC_8_8_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i26_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i26_LC_8_8_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i26_LC_8_8_4  (
            .in0(N__24099),
            .in1(N__34962),
            .in2(N__34826),
            .in3(N__35672),
            .lcout(cmd_33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i11_LC_8_8_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i11_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i11_LC_8_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i11_LC_8_8_5  (
            .in0(N__35477),
            .in1(N__34592),
            .in2(_gnd_net_),
            .in3(N__24283),
            .lcout(bwd_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i28_LC_8_8_6 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i28_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i28_LC_8_8_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i28_LC_8_8_6  (
            .in0(N__24371),
            .in1(N__34963),
            .in2(N__28176),
            .in3(N__34803),
            .lcout(cmd_35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i21_LC_8_8_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i21_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i21_LC_8_8_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i21_LC_8_8_7  (
            .in0(N__24152),
            .in1(_gnd_net_),
            .in2(N__34119),
            .in3(N__24117),
            .lcout(configRegister_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i4_LC_8_9_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i4_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i4_LC_8_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i4_LC_8_9_0  (
            .in0(N__29114),
            .in1(N__26752),
            .in2(_gnd_net_),
            .in3(N__35510),
            .lcout(bwd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i2_LC_8_9_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i2_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i2_LC_8_9_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i2_LC_8_9_1  (
            .in0(N__35509),
            .in1(_gnd_net_),
            .in2(N__29691),
            .in3(N__29932),
            .lcout(bwd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i29_LC_8_9_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i29_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i29_LC_8_9_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i29_LC_8_9_2  (
            .in0(N__34799),
            .in1(N__35053),
            .in2(N__24395),
            .in3(N__24366),
            .lcout(cmd_36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i9_LC_8_9_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i9_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i9_LC_8_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i9_LC_8_9_3  (
            .in0(N__35514),
            .in1(N__24100),
            .in2(_gnd_net_),
            .in3(N__24199),
            .lcout(fwd_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i13_LC_8_9_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i13_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i13_LC_8_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i13_LC_8_9_4  (
            .in0(N__24391),
            .in1(N__35512),
            .in2(_gnd_net_),
            .in3(N__24212),
            .lcout(fwd_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i1_LC_8_9_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i1_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i1_LC_8_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i1_LC_8_9_5  (
            .in0(N__35513),
            .in1(N__29540),
            .in2(_gnd_net_),
            .in3(N__24484),
            .lcout(fwd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i12_LC_8_9_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i12_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i12_LC_8_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i12_LC_8_9_6  (
            .in0(N__24502),
            .in1(N__24367),
            .in2(_gnd_net_),
            .in3(N__35511),
            .lcout(fwd_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i7_LC_8_9_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i7_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i7_LC_8_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i7_LC_8_9_7  (
            .in0(N__35831),
            .in1(N__24346),
            .in2(_gnd_net_),
            .in3(N__34423),
            .lcout(configRegister_6_adj_1354),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i5_LC_8_10_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i5_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i5_LC_8_10_0 .LUT_INIT=16'b0110011001011010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i5_LC_8_10_0  (
            .in0(N__24335),
            .in1(N__24317),
            .in2(N__25514),
            .in3(N__30332),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37547),
            .ce(),
            .sr(N__24296));
    defparam \Inst_core.Inst_controller.i2_4_lut_adj_60_LC_8_10_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i2_4_lut_adj_60_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i2_4_lut_adj_60_LC_8_10_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_controller.i2_4_lut_adj_60_LC_8_10_1  (
            .in0(N__37772),
            .in1(N__24284),
            .in2(N__24269),
            .in3(N__36929),
            .lcout(\Inst_core.Inst_controller.n18_adj_990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i6_4_lut_LC_8_10_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i6_4_lut_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i6_4_lut_LC_8_10_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_controller.i6_4_lut_LC_8_10_2  (
            .in0(N__24250),
            .in1(N__37078),
            .in2(N__26486),
            .in3(N__37771),
            .lcout(),
            .ltout(\Inst_core.Inst_controller.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i9_4_lut_LC_8_10_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i9_4_lut_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i9_4_lut_LC_8_10_3 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \Inst_core.Inst_controller.i9_4_lut_LC_8_10_3  (
            .in0(N__24235),
            .in1(N__37051),
            .in2(N__24221),
            .in3(N__24422),
            .lcout(\Inst_core.Inst_controller.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i3_4_lut_LC_8_10_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i3_4_lut_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i3_4_lut_LC_8_10_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_controller.i3_4_lut_LC_8_10_4  (
            .in0(N__24211),
            .in1(N__36901),
            .in2(N__24200),
            .in3(N__37724),
            .lcout(\Inst_core.Inst_controller.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i4_LC_8_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i4_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i4_LC_8_11_0 .LUT_INIT=16'b0010110101111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i4_LC_8_11_0  (
            .in0(N__30358),
            .in1(N__24587),
            .in2(N__24560),
            .in3(N__28085),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37559),
            .ce(),
            .sr(N__24539));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_adj_71_LC_8_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_adj_71_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_adj_71_LC_8_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3_4_lut_adj_71_LC_8_11_1  (
            .in0(N__24527),
            .in1(N__30233),
            .in2(N__24521),
            .in3(N__24509),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i1_4_lut_LC_8_11_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1_4_lut_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1_4_lut_LC_8_11_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_controller.i1_4_lut_LC_8_11_2  (
            .in0(N__24503),
            .in1(N__36211),
            .in2(N__24488),
            .in3(N__37747),
            .lcout(\Inst_core.Inst_controller.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i4_4_lut_adj_59_LC_8_11_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i4_4_lut_adj_59_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i4_4_lut_adj_59_LC_8_11_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \Inst_core.Inst_controller.i4_4_lut_adj_59_LC_8_11_3  (
            .in0(N__37748),
            .in1(N__24464),
            .in2(N__35240),
            .in3(N__37796),
            .lcout(\Inst_core.Inst_controller.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i8_4_lut_LC_8_11_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i8_4_lut_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i8_4_lut_LC_8_11_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \Inst_core.Inst_controller.i8_4_lut_LC_8_11_4  (
            .in0(N__34142),
            .in1(N__36953),
            .in2(N__36215),
            .in3(N__27076),
            .lcout(\Inst_core.Inst_controller.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i2_4_lut_LC_8_11_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i2_4_lut_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i2_4_lut_LC_8_11_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \Inst_core.Inst_controller.i2_4_lut_LC_8_11_5  (
            .in0(N__36952),
            .in1(N__27064),
            .in2(N__28985),
            .in3(N__37795),
            .lcout(\Inst_core.Inst_controller.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.counter_17__I_0_43_i11_2_lut_LC_8_11_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.counter_17__I_0_43_i11_2_lut_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.counter_17__I_0_43_i11_2_lut_LC_8_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Inst_core.Inst_controller.counter_17__I_0_43_i11_2_lut_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__24443),
            .in2(_gnd_net_),
            .in3(N__36928),
            .lcout(\Inst_core.Inst_controller.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register_80_LC_8_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register_80_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register_80_LC_8_12_0 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register_80_LC_8_12_0  (
            .in0(N__24416),
            .in1(N__24401),
            .in2(_gnd_net_),
            .in3(N__26362),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.match32Register ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i1_LC_8_12_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i1_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i1_LC_8_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i1_LC_8_12_1  (
            .in0(N__27051),
            .in1(N__34257),
            .in2(_gnd_net_),
            .in3(N__27476),
            .lcout(maskRegister_1_adj_1327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i21_LC_8_12_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i21_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i21_LC_8_12_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i21_LC_8_12_2  (
            .in0(N__24686),
            .in1(N__31168),
            .in2(_gnd_net_),
            .in3(N__25027),
            .lcout(divider_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i0_LC_8_12_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i0_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i0_LC_8_12_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i0_LC_8_12_3  (
            .in0(N__31166),
            .in1(N__24635),
            .in2(N__31788),
            .in3(N__31953),
            .lcout(memoryOut_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i4_LC_8_12_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i4_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i4_LC_8_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i4_LC_8_12_4  (
            .in0(N__29494),
            .in1(N__24607),
            .in2(_gnd_net_),
            .in3(N__29132),
            .lcout(valueRegister_4_adj_1332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3597_1_lut_LC_8_12_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3597_1_lut_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3597_1_lut_LC_8_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3597_1_lut_LC_8_12_5  (
            .in0(N__26980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i1_LC_8_12_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i1_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i1_LC_8_12_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i1_LC_8_12_6  (
            .in0(N__34258),
            .in1(_gnd_net_),
            .in2(N__29495),
            .in3(N__25066),
            .lcout(valueRegister_1_adj_1335),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.sample_i0_i1_LC_8_12_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.sample_i0_i1_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.sample_i0_i1_LC_8_12_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Inst_core.Inst_sampler.sample_i0_i1_LC_8_12_7  (
            .in0(N__31167),
            .in1(N__33608),
            .in2(N__24629),
            .in3(N__31954),
            .lcout(memoryOut_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i4_LC_8_13_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i4_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i4_LC_8_13_0 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i4_LC_8_13_0  (
            .in0(N__25145),
            .in1(N__35606),
            .in2(N__24614),
            .in3(N__28072),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37586),
            .ce(),
            .sr(N__24596));
    defparam \Inst_core.Inst_sampler.i7_4_lut_LC_8_13_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7_4_lut_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7_4_lut_LC_8_13_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i7_4_lut_LC_8_13_1  (
            .in0(N__25023),
            .in1(N__27850),
            .in2(N__29971),
            .in3(N__27805),
            .lcout(),
            .ltout(\Inst_core.Inst_sampler.n31_adj_995_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i20_4_lut_LC_8_13_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i20_4_lut_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i20_4_lut_LC_8_13_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_sampler.i20_4_lut_LC_8_13_2  (
            .in0(N__24731),
            .in1(N__27332),
            .in2(N__24590),
            .in3(N__24848),
            .lcout(\Inst_core.Inst_sampler.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i5_4_lut_LC_8_13_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i5_4_lut_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i5_4_lut_LC_8_13_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i5_4_lut_LC_8_13_3  (
            .in0(N__24895),
            .in1(N__27525),
            .in2(N__24872),
            .in3(N__27701),
            .lcout(\Inst_core.Inst_sampler.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_adj_72_LC_8_13_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_adj_72_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_adj_72_LC_8_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_adj_72_LC_8_13_4  (
            .in0(N__27383),
            .in1(N__24842),
            .in2(N__24812),
            .in3(N__24833),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7_adj_996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i5_LC_8_14_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i5_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i5_LC_8_14_0 .LUT_INIT=16'b0010011111011000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i5_LC_8_14_0  (
            .in0(N__35601),
            .in1(N__25124),
            .in2(N__25511),
            .in3(N__24827),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37597),
            .ce(),
            .sr(N__25883));
    defparam \Inst_core.Inst_sampler.i4_4_lut_LC_8_14_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i4_4_lut_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i4_4_lut_LC_8_14_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i4_4_lut_LC_8_14_1  (
            .in0(N__24801),
            .in1(N__27648),
            .in2(N__24778),
            .in3(N__27612),
            .lcout(\Inst_core.Inst_sampler.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7236_4_lut_LC_8_14_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7236_4_lut_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7236_4_lut_LC_8_14_2 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_sampler.i7236_4_lut_LC_8_14_2  (
            .in0(N__24802),
            .in1(N__27631),
            .in2(N__24785),
            .in3(N__31548),
            .lcout(\Inst_core.Inst_sampler.n8604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7230_4_lut_LC_8_14_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7230_4_lut_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7230_4_lut_LC_8_14_3 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_sampler.i7230_4_lut_LC_8_14_3  (
            .in0(N__24748),
            .in1(N__27613),
            .in2(N__29975),
            .in3(N__30617),
            .lcout(\Inst_core.Inst_sampler.n8598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i8_4_lut_LC_8_14_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i8_4_lut_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i8_4_lut_LC_8_14_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i8_4_lut_LC_8_14_4  (
            .in0(N__24747),
            .in1(N__27630),
            .in2(N__24724),
            .in3(N__27592),
            .lcout(\Inst_core.Inst_sampler.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7228_4_lut_LC_8_14_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7228_4_lut_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7228_4_lut_LC_8_14_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i7228_4_lut_LC_8_14_5  (
            .in0(N__27299),
            .in1(N__27649),
            .in2(N__24725),
            .in3(N__27699),
            .lcout(),
            .ltout(\Inst_core.Inst_sampler.n8596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7300_4_lut_LC_8_14_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7300_4_lut_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7300_4_lut_LC_8_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_sampler.i7300_4_lut_LC_8_14_6  (
            .in0(N__27215),
            .in1(N__27326),
            .in2(N__24695),
            .in3(N__24692),
            .lcout(\Inst_core.Inst_sampler.n8669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i1_LC_8_15_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i1_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i1_LC_8_15_0 .LUT_INIT=16'b0110010101101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i1_LC_8_15_0  (
            .in0(N__25070),
            .in1(N__24914),
            .in2(N__35611),
            .in3(N__33633),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37606),
            .ce(),
            .sr(N__27464));
    defparam \Inst_core.Inst_sampler.i11_4_lut_LC_8_15_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i11_4_lut_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i11_4_lut_LC_8_15_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i11_4_lut_LC_8_15_1  (
            .in0(N__25055),
            .in1(N__27876),
            .in2(N__27248),
            .in3(N__27822),
            .lcout(\Inst_core.Inst_sampler.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7232_4_lut_LC_8_15_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7232_4_lut_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7232_4_lut_LC_8_15_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \Inst_core.Inst_sampler.i7232_4_lut_LC_8_15_2  (
            .in0(N__27823),
            .in1(N__27362),
            .in2(N__25031),
            .in3(N__30501),
            .lcout(),
            .ltout(\Inst_core.Inst_sampler.n8600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7302_4_lut_LC_8_15_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7302_4_lut_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7302_4_lut_LC_8_15_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_sampler.i7302_4_lut_LC_8_15_3  (
            .in0(N__25007),
            .in1(N__24998),
            .in2(N__24989),
            .in3(N__24986),
            .lcout(\Inst_core.Inst_sampler.n8671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i0_LC_8_16_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i0_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i0_LC_8_16_0 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i0_LC_8_16_0  (
            .in0(N__26390),
            .in1(N__24937),
            .in2(N__24980),
            .in3(N__24956),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i1_LC_8_16_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i1_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i1_LC_8_16_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i1_LC_8_16_1  (
            .in0(N__24938),
            .in1(N__32190),
            .in2(_gnd_net_),
            .in3(N__26383),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i2_LC_8_16_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i2_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i2_LC_8_16_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i2_LC_8_16_2  (
            .in0(N__26384),
            .in1(_gnd_net_),
            .in2(N__32197),
            .in3(N__24912),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i3_LC_8_16_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i3_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i3_LC_8_16_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i3_LC_8_16_3  (
            .in0(N__24913),
            .in1(N__30816),
            .in2(_gnd_net_),
            .in3(N__26385),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i4_LC_8_16_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i4_LC_8_16_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i4_LC_8_16_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i4_LC_8_16_4  (
            .in0(N__26386),
            .in1(_gnd_net_),
            .in2(N__30823),
            .in3(N__31617),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i5_LC_8_16_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i5_LC_8_16_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i5_LC_8_16_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i5_LC_8_16_5  (
            .in0(N__31618),
            .in1(N__25137),
            .in2(_gnd_net_),
            .in3(N__26387),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i6_LC_8_16_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i6_LC_8_16_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i6_LC_8_16_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i6_LC_8_16_6  (
            .in0(N__26388),
            .in1(_gnd_net_),
            .in2(N__25144),
            .in3(N__25119),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i7_LC_8_16_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i7_LC_8_16_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i7_LC_8_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_i0_i7_LC_8_16_7  (
            .in0(N__25120),
            .in1(N__27415),
            .in2(_gnd_net_),
            .in3(N__26389),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.shiftRegister_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7564_4_lut_LC_9_1_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7564_4_lut_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7564_4_lut_LC_9_1_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i7564_4_lut_LC_9_1_0  (
            .in0(N__25365),
            .in1(N__27723),
            .in2(N__36657),
            .in3(N__25746),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n8844_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.run_83_LC_9_1_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.run_83_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.run_83_LC_9_1_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.run_83_LC_9_1_1  (
            .in0(N__36859),
            .in1(_gnd_net_),
            .in2(N__25091),
            .in3(N__32524),
            .lcout(\Inst_core.Inst_trigger.stageRun_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37616),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.run_83_LC_9_1_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.run_83_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.run_83_LC_9_1_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.run_83_LC_9_1_2  (
            .in0(N__32440),
            .in1(N__36860),
            .in2(_gnd_net_),
            .in3(N__32555),
            .lcout(\Inst_core.Inst_trigger.stageRun_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37616),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.run_83_LC_9_1_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.run_83_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.run_83_LC_9_1_3 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.run_83_LC_9_1_3  (
            .in0(N__25185),
            .in1(_gnd_net_),
            .in2(N__36874),
            .in3(N__25088),
            .lcout(\Inst_core.stageRun_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37616),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7644_4_lut_LC_9_1_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7644_4_lut_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7644_4_lut_LC_9_1_4 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i7644_4_lut_LC_9_1_4  (
            .in0(N__25366),
            .in1(N__25745),
            .in2(N__36656),
            .in3(N__36858),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n8622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7667_1_lut_2_lut_3_lut_LC_9_1_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7667_1_lut_2_lut_3_lut_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i7667_1_lut_2_lut_3_lut_LC_9_1_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i7667_1_lut_2_lut_3_lut_LC_9_1_5  (
            .in0(N__25743),
            .in1(N__36625),
            .in2(_gnd_net_),
            .in3(N__25363),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n9052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i25_LC_9_1_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i25_LC_9_1_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i25_LC_9_1_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i25_LC_9_1_6  (
            .in0(N__26106),
            .in1(N__28199),
            .in2(_gnd_net_),
            .in3(N__27724),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister_27_adj_997 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37616),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i890_2_lut_3_lut_LC_9_1_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i890_2_lut_3_lut_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i890_2_lut_3_lut_LC_9_1_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i890_2_lut_3_lut_LC_9_1_7  (
            .in0(N__25744),
            .in1(N__36626),
            .in2(_gnd_net_),
            .in3(N__25364),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n1765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i199_2_lut_3_lut_LC_9_2_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i199_2_lut_3_lut_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i199_2_lut_3_lut_LC_9_2_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i199_2_lut_3_lut_LC_9_2_0  (
            .in0(N__25204),
            .in1(N__26188),
            .in2(_gnd_net_),
            .in3(N__28879),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n667 ),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n667_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i3_LC_9_2_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i3_LC_9_2_1 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i3_LC_9_2_1 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i3_LC_9_2_1  (
            .in0(N__36663),
            .in1(N__25186),
            .in2(N__25235),
            .in3(N__25232),
            .lcout(\Inst_core.state_1_adj_1134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37609),
            .ce(),
            .sr(N__36865));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i44_2_lut_LC_9_2_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i44_2_lut_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i44_2_lut_LC_9_2_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i44_2_lut_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__26189),
            .in2(_gnd_net_),
            .in3(N__28880),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i2_LC_9_2_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i2_LC_9_2_3 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i2_LC_9_2_3 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i2_LC_9_2_3  (
            .in0(N__25154),
            .in1(N__25934),
            .in2(N__25208),
            .in3(N__25205),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37609),
            .ce(),
            .sr(N__36865));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i3_LC_9_2_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i3_LC_9_2_4 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i3_LC_9_2_4 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i3_LC_9_2_4  (
            .in0(N__28326),
            .in1(N__32957),
            .in2(N__27911),
            .in3(N__36664),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37609),
            .ce(),
            .sr(N__36865));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i1_LC_9_2_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i1_LC_9_2_5 .SEQ_MODE=4'b1011;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i1_LC_9_2_5 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.state_FSM_i1_LC_9_2_5  (
            .in0(N__25153),
            .in1(N__25196),
            .in2(N__25190),
            .in3(N__25935),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37609),
            .ce(),
            .sr(N__36865));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i1_LC_9_2_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i1_LC_9_2_6 .SEQ_MODE=4'b1011;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i1_LC_9_2_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i1_LC_9_2_6  (
            .in0(N__25932),
            .in1(N__25399),
            .in2(_gnd_net_),
            .in3(N__28358),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37609),
            .ce(),
            .sr(N__36865));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i2_LC_9_2_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i2_LC_9_2_7 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i2_LC_9_2_7 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.state_FSM_i2_LC_9_2_7  (
            .in0(N__25841),
            .in1(N__25933),
            .in2(N__25403),
            .in3(N__25831),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37609),
            .ce(),
            .sr(N__36865));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_LC_9_3_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_LC_9_3_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__25739),
            .in2(_gnd_net_),
            .in3(N__25361),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i1_LC_9_3_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i1_LC_9_3_1 .SEQ_MODE=4'b1011;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i1_LC_9_3_1 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i1_LC_9_3_1  (
            .in0(N__25937),
            .in1(N__36646),
            .in2(N__25391),
            .in3(N__25375),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(N__36864));
    defparam \Inst_core.Inst_sampler.i1_2_lut_LC_9_3_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i1_2_lut_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i1_2_lut_LC_9_3_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Inst_core.Inst_sampler.i1_2_lut_LC_9_3_2  (
            .in0(N__36645),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32433),
            .lcout(),
            .ltout(\Inst_core.n8515_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i1_LC_9_3_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i1_LC_9_3_3 .SEQ_MODE=4'b1011;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i1_LC_9_3_3 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i1_LC_9_3_3  (
            .in0(N__25939),
            .in1(N__25384),
            .in2(N__25388),
            .in3(N__33268),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(N__36864));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i2_LC_9_3_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i2_LC_9_3_4 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i2_LC_9_3_4 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i2_LC_9_3_4  (
            .in0(N__25385),
            .in1(N__25936),
            .in2(N__28573),
            .in3(N__28589),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(N__36864));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i2_LC_9_3_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i2_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i2_LC_9_3_5 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i2_LC_9_3_5  (
            .in0(N__25938),
            .in1(N__25376),
            .in2(N__25775),
            .in3(N__25787),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(N__36864));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i3_LC_9_3_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i3_LC_9_3_6 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i3_LC_9_3_6 .LUT_INIT=16'b1111111110001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.state_FSM_i3_LC_9_3_6  (
            .in0(N__33269),
            .in1(N__32434),
            .in2(N__36662),
            .in3(N__32474),
            .lcout(\Inst_core.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(N__36864));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i3_LC_9_3_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i3_LC_9_3_7 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i3_LC_9_3_7 .LUT_INIT=16'b1111111110110000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.state_FSM_i3_LC_9_3_7  (
            .in0(N__25362),
            .in1(N__36647),
            .in2(N__25748),
            .in3(N__25757),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(N__36864));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register_80_LC_9_4_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register_80_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register_80_LC_9_4_0 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register_80_LC_9_4_0  (
            .in0(N__32675),
            .in1(N__27926),
            .in2(_gnd_net_),
            .in3(N__26382),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.match32Register ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i6_LC_9_4_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i6_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i6_LC_9_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i6_LC_9_4_1  (
            .in0(N__29252),
            .in1(N__28549),
            .in2(_gnd_net_),
            .in3(N__31383),
            .lcout(configRegister_5_adj_1315),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i10_LC_9_4_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i10_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i10_LC_9_4_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i10_LC_9_4_2  (
            .in0(N__25599),
            .in1(N__31031),
            .in2(_gnd_net_),
            .in3(N__27294),
            .lcout(divider_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i4_LC_9_4_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i4_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i4_LC_9_4_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i4_LC_9_4_3  (
            .in0(N__29251),
            .in1(N__28234),
            .in2(_gnd_net_),
            .in3(N__26725),
            .lcout(configRegister_3_adj_1317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i14_LC_9_4_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i14_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i14_LC_9_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i14_LC_9_4_4  (
            .in0(N__35858),
            .in1(N__29355),
            .in2(_gnd_net_),
            .in3(N__25558),
            .lcout(configRegister_13_adj_1347),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i15_LC_9_4_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i15_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i15_LC_9_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i15_LC_9_4_5  (
            .in0(N__26137),
            .in1(N__30115),
            .in2(_gnd_net_),
            .in3(N__25543),
            .lcout(configRegister_14_adj_1386),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i7_LC_9_4_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i7_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i7_LC_9_4_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i7_LC_9_4_6  (
            .in0(N__34433),
            .in1(N__29253),
            .in2(_gnd_net_),
            .in3(N__28531),
            .lcout(configRegister_6_adj_1314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i3_LC_9_4_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i3_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i3_LC_9_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i3_LC_9_4_7  (
            .in0(N__29250),
            .in1(N__28255),
            .in2(_gnd_net_),
            .in3(N__29675),
            .lcout(configRegister_2_adj_1318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37589),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i5_LC_9_5_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i5_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i5_LC_9_5_0 .LUT_INIT=16'b0110011001011010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i5_LC_9_5_0  (
            .in0(N__26177),
            .in1(N__25532),
            .in2(N__25507),
            .in3(N__33551),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37576),
            .ce(),
            .sr(N__25625));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_2_lut_LC_9_5_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_2_lut_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_2_lut_LC_9_5_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_2_lut_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__26612),
            .in2(_gnd_net_),
            .in3(N__28956),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i44_4_lut_LC_9_5_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i44_4_lut_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i44_4_lut_LC_9_5_2 .LUT_INIT=16'b0100110100000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i44_4_lut_LC_9_5_2  (
            .in0(N__25673),
            .in1(N__28910),
            .in2(N__25856),
            .in3(N__25853),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n100 ),
            .ltout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i166_2_lut_LC_9_5_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i166_2_lut_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i166_2_lut_LC_9_5_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i166_2_lut_LC_9_5_3  (
            .in0(N__25832),
            .in1(_gnd_net_),
            .in2(N__25817),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_74_LC_9_5_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_74_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_74_LC_9_5_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_74_LC_9_5_4  (
            .in0(N__28957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25970),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i44_4_lut_LC_9_5_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i44_4_lut_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i44_4_lut_LC_9_5_5 .LUT_INIT=16'b0000100010001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i44_4_lut_LC_9_5_5  (
            .in0(N__28911),
            .in1(N__25814),
            .in2(N__25808),
            .in3(N__25805),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n100 ),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i232_2_lut_LC_9_5_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i232_2_lut_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i232_2_lut_LC_9_5_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i232_2_lut_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25778),
            .in3(N__25774),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n770 ),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n770_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_4_lut_adj_75_LC_9_5_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_4_lut_adj_75_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_4_lut_adj_75_LC_9_5_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_4_lut_adj_75_LC_9_5_7  (
            .in0(N__25747),
            .in1(N__36808),
            .in2(N__25709),
            .in3(N__25706),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4076 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i18_LC_9_6_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i18_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i18_LC_9_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i18_LC_9_6_0  (
            .in0(N__29318),
            .in1(N__29548),
            .in2(_gnd_net_),
            .in3(N__25672),
            .lcout(configRegister_17_adj_1303),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i5_LC_9_6_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i5_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i5_LC_9_6_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i5_LC_9_6_1  (
            .in0(N__29122),
            .in1(N__35835),
            .in2(_gnd_net_),
            .in3(N__25651),
            .lcout(configRegister_4_adj_1356),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3605_1_lut_LC_9_6_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3605_1_lut_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3605_1_lut_LC_9_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3605_1_lut_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25640),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i10_LC_9_6_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i10_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i10_LC_9_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i10_LC_9_6_3  (
            .in0(N__34096),
            .in1(N__33109),
            .in2(_gnd_net_),
            .in3(N__26595),
            .lcout(configRegister_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i10_LC_9_6_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i10_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i10_LC_9_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i10_LC_9_6_4  (
            .in0(N__26594),
            .in1(N__29320),
            .in2(_gnd_net_),
            .in3(N__28462),
            .lcout(configRegister_9_adj_1311),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i13_LC_9_6_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i13_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i13_LC_9_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i13_LC_9_6_5  (
            .in0(N__35289),
            .in1(N__35834),
            .in2(_gnd_net_),
            .in3(N__25951),
            .lcout(configRegister_12_adj_1348),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i5_LC_9_6_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i5_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i5_LC_9_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i5_LC_9_6_6  (
            .in0(N__29319),
            .in1(N__28213),
            .in2(_gnd_net_),
            .in3(N__29123),
            .lcout(configRegister_4_adj_1316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i15_LC_9_6_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i15_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i15_LC_9_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i15_LC_9_6_7  (
            .in0(N__34097),
            .in1(N__30100),
            .in2(_gnd_net_),
            .in3(N__33814),
            .lcout(configRegister_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.levelReg_927__i1_LC_9_7_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.levelReg_927__i1_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.levelReg_927__i1_LC_9_7_0 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \Inst_core.Inst_trigger.levelReg_927__i1_LC_9_7_0  (
            .in0(N__28955),
            .in1(_gnd_net_),
            .in2(N__33368),
            .in3(N__28909),
            .lcout(\Inst_core.Inst_trigger.levelReg_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37549),
            .ce(),
            .sr(N__25940));
    defparam \Inst_core.Inst_trigger.levelReg_927__i0_LC_9_7_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.levelReg_927__i0_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_trigger.levelReg_927__i0_LC_9_7_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Inst_core.Inst_trigger.levelReg_927__i0_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__33364),
            .in2(_gnd_net_),
            .in3(N__28954),
            .lcout(\Inst_core.Inst_trigger.levelReg_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37549),
            .ce(),
            .sr(N__25940));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3598_1_lut_LC_9_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3598_1_lut_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3598_1_lut_LC_9_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3598_1_lut_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25894),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3599_1_lut_LC_9_7_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3599_1_lut_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3599_1_lut_LC_9_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3599_1_lut_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25867),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3600_1_lut_LC_9_7_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3600_1_lut_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3600_1_lut_LC_9_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3600_1_lut_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26471),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3486_1_lut_LC_9_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3486_1_lut_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3486_1_lut_LC_9_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3486_1_lut_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26437),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3601_1_lut_LC_9_7_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3601_1_lut_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3601_1_lut_LC_9_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3601_1_lut_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26425),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3602_1_lut_LC_9_7_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3602_1_lut_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3602_1_lut_LC_9_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3602_1_lut_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26413),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n4761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register_80_LC_9_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register_80_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register_80_LC_9_8_0 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register_80_LC_9_8_0  (
            .in0(N__32123),
            .in1(N__26402),
            .in2(_gnd_net_),
            .in3(N__26381),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.match32Register ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i5_LC_9_8_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i5_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i5_LC_9_8_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i5_LC_9_8_1  (
            .in0(N__31332),
            .in1(N__36103),
            .in2(_gnd_net_),
            .in3(N__26173),
            .lcout(valueRegister_5_adj_1371),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i0_LC_9_8_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i0_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i0_LC_9_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i0_LC_9_8_2  (
            .in0(N__30205),
            .in1(N__36175),
            .in2(_gnd_net_),
            .in3(N__35466),
            .lcout(fwd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i14_LC_9_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i14_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i14_LC_9_8_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i14_LC_9_8_3  (
            .in0(N__29394),
            .in1(N__26144),
            .in2(_gnd_net_),
            .in3(N__26155),
            .lcout(configRegister_13_adj_1387),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i17_LC_9_8_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i17_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i17_LC_9_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.configRegister__i17_LC_9_8_4  (
            .in0(N__26143),
            .in1(N__36177),
            .in2(_gnd_net_),
            .in3(N__25969),
            .lcout(configRegister_16_adj_1384),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i17_LC_9_8_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i17_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i17_LC_9_8_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i17_LC_9_8_5  (
            .in0(N__36176),
            .in1(N__29325),
            .in2(_gnd_net_),
            .in3(N__26611),
            .lcout(configRegister_16_adj_1304),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i9_LC_9_8_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i9_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i9_LC_9_8_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i9_LC_9_8_7  (
            .in0(N__35465),
            .in1(N__26587),
            .in2(_gnd_net_),
            .in3(N__26887),
            .lcout(bwd_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i13_LC_9_9_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i13_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i13_LC_9_9_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i13_LC_9_9_0  (
            .in0(N__35270),
            .in1(N__34821),
            .in2(N__29399),
            .in3(N__35055),
            .lcout(cmd_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i20_LC_9_9_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i20_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i20_LC_9_9_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i20_LC_9_9_1  (
            .in0(N__35054),
            .in1(N__26540),
            .in2(N__34842),
            .in3(N__29988),
            .lcout(cmd_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i6_LC_9_9_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i6_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i6_LC_9_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i6_LC_9_9_2  (
            .in0(N__35516),
            .in1(N__34428),
            .in2(_gnd_net_),
            .in3(N__26801),
            .lcout(bwd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i3_LC_9_9_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i3_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i3_LC_9_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i3_LC_9_9_3  (
            .in0(N__26729),
            .in1(N__29475),
            .in2(_gnd_net_),
            .in3(N__31594),
            .lcout(valueRegister_3_adj_1333),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i3_LC_9_9_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i3_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i3_LC_9_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i3_LC_9_9_4  (
            .in0(N__27049),
            .in1(N__26728),
            .in2(_gnd_net_),
            .in3(N__27436),
            .lcout(maskRegister_3_adj_1325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i3_LC_9_9_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i3_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i3_LC_9_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i3_LC_9_9_5  (
            .in0(N__26727),
            .in1(N__34521),
            .in2(_gnd_net_),
            .in3(N__26842),
            .lcout(valueRegister_3_adj_1293),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i3_LC_9_9_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i3_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i3_LC_9_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i3_LC_9_9_6  (
            .in0(N__35515),
            .in1(N__26726),
            .in2(_gnd_net_),
            .in3(N__26765),
            .lcout(bwd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i3_LC_9_9_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i3_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i3_LC_9_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i3_LC_9_9_7  (
            .in0(N__35517),
            .in1(N__29989),
            .in2(_gnd_net_),
            .in3(N__26485),
            .lcout(fwd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i6_4_lut_adj_58_LC_9_10_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i6_4_lut_adj_58_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i6_4_lut_adj_58_LC_9_10_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_controller.i6_4_lut_adj_58_LC_9_10_0  (
            .in0(N__26888),
            .in1(N__37664),
            .in2(N__28832),
            .in3(N__36902),
            .lcout(),
            .ltout(\Inst_core.Inst_controller.n22_adj_988_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i14_4_lut_LC_9_10_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i14_4_lut_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i14_4_lut_LC_9_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_controller.i14_4_lut_LC_9_10_1  (
            .in0(N__26873),
            .in1(N__26771),
            .in2(N__26867),
            .in3(N__26738),
            .lcout(\Inst_core.Inst_controller.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i3_LC_9_10_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i3_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i3_LC_9_10_2 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i3_LC_9_10_2  (
            .in0(N__26864),
            .in1(N__26843),
            .in2(N__30346),
            .in3(N__32351),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37561),
            .ce(),
            .sr(N__26813));
    defparam \Inst_core.Inst_controller.i7_4_lut_LC_9_10_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i7_4_lut_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i7_4_lut_LC_9_10_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_controller.i7_4_lut_LC_9_10_3  (
            .in0(N__26800),
            .in1(N__37024),
            .in2(N__26789),
            .in3(N__36988),
            .lcout(\Inst_core.Inst_controller.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i5_4_lut_LC_9_10_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i5_4_lut_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i5_4_lut_LC_9_10_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \Inst_core.Inst_controller.i5_4_lut_LC_9_10_4  (
            .in0(N__37052),
            .in1(N__26764),
            .in2(N__26753),
            .in3(N__37079),
            .lcout(\Inst_core.Inst_controller.n21_adj_989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i2_LC_9_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i2_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i2_LC_9_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i2_LC_9_11_0  (
            .in0(N__31112),
            .in1(N__29713),
            .in2(_gnd_net_),
            .in3(N__27315),
            .lcout(divider_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i18_LC_9_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i18_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i18_LC_9_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i18_LC_9_11_1  (
            .in0(N__30035),
            .in1(N__31114),
            .in2(_gnd_net_),
            .in3(N__30579),
            .lcout(divider_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i3_LC_9_11_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i3_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i3_LC_9_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i3_LC_9_11_2  (
            .in0(N__31113),
            .in1(N__26731),
            .in2(_gnd_net_),
            .in3(N__31683),
            .lcout(divider_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i2_LC_9_11_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i2_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i2_LC_9_11_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i2_LC_9_11_3  (
            .in0(N__29711),
            .in1(N__27042),
            .in2(_gnd_net_),
            .in3(N__27449),
            .lcout(maskRegister_2_adj_1326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i7_LC_9_11_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i7_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i7_LC_9_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i7_LC_9_11_4  (
            .in0(N__35518),
            .in1(N__27207),
            .in2(_gnd_net_),
            .in3(N__27077),
            .lcout(bwd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i2_LC_9_11_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i2_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i2_LC_9_11_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i2_LC_9_11_5  (
            .in0(N__29712),
            .in1(N__29490),
            .in2(_gnd_net_),
            .in3(N__30838),
            .lcout(valueRegister_2_adj_1334),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i10_LC_9_11_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i10_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i10_LC_9_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i10_LC_9_11_6  (
            .in0(N__35519),
            .in1(N__35680),
            .in2(_gnd_net_),
            .in3(N__27065),
            .lcout(fwd_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i4_LC_9_11_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i4_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i4_LC_9_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.maskRegister_i0_i4_LC_9_11_7  (
            .in0(N__27043),
            .in1(N__29129),
            .in2(_gnd_net_),
            .in3(N__26981),
            .lcout(maskRegister_4_adj_1324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.result_i7_LC_9_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i7_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.result_i7_LC_9_12_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.result_i7_LC_9_12_0  (
            .in0(N__26962),
            .in1(N__31472),
            .in2(_gnd_net_),
            .in3(N__31436),
            .lcout(\Inst_core.Inst_sync.filteredInput_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37588),
            .ce(),
            .sr(N__26948));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3593_1_lut_LC_9_12_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3593_1_lut_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3593_1_lut_LC_9_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3593_1_lut_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26936),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7670_1_lut_LC_9_12_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7670_1_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7670_1_lut_LC_9_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i7670_1_lut_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28769),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n9055 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3484_1_lut_LC_9_12_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3484_1_lut_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3484_1_lut_LC_9_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3484_1_lut_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26903),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3594_1_lut_LC_9_12_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3594_1_lut_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3594_1_lut_LC_9_12_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3594_1_lut_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__27475),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3595_1_lut_LC_9_12_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3595_1_lut_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3595_1_lut_LC_9_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3595_1_lut_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27448),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3596_1_lut_LC_9_12_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3596_1_lut_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3596_1_lut_LC_9_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3596_1_lut_LC_9_12_6  (
            .in0(N__27437),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n4755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i6_LC_9_13_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i6_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i6_LC_9_13_0 .LUT_INIT=16'b0011010111001010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i6_LC_9_13_0  (
            .in0(N__30452),
            .in1(N__27422),
            .in2(N__35600),
            .in3(N__27404),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37599),
            .ce(),
            .sr(N__27377));
    defparam \Inst_core.Inst_sampler.i6_4_lut_LC_9_13_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i6_4_lut_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i6_4_lut_LC_9_13_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_sampler.i6_4_lut_LC_9_13_1  (
            .in0(N__30699),
            .in1(N__27316),
            .in2(N__27361),
            .in3(N__27552),
            .lcout(\Inst_core.Inst_sampler.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7224_4_lut_LC_9_13_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7224_4_lut_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7224_4_lut_LC_9_13_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i7224_4_lut_LC_9_13_2  (
            .in0(N__27274),
            .in1(N__27553),
            .in2(N__32108),
            .in3(N__27526),
            .lcout(\Inst_core.Inst_sampler.n8592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7238_4_lut_LC_9_13_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7238_4_lut_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7238_4_lut_LC_9_13_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \Inst_core.Inst_sampler.i7238_4_lut_LC_9_13_3  (
            .in0(N__30583),
            .in1(N__30555),
            .in2(N__27887),
            .in3(N__27317),
            .lcout(\Inst_core.Inst_sampler.n8606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i9_4_lut_LC_9_13_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i9_4_lut_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i9_4_lut_LC_9_13_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i9_4_lut_LC_9_13_4  (
            .in0(N__27295),
            .in1(N__27502),
            .in2(N__27275),
            .in3(N__27676),
            .lcout(\Inst_core.Inst_sampler.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7220_4_lut_LC_9_13_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7220_4_lut_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7220_4_lut_LC_9_13_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i7220_4_lut_LC_9_13_5  (
            .in0(N__27677),
            .in1(N__27247),
            .in2(N__27596),
            .in3(N__30785),
            .lcout(\Inst_core.Inst_sampler.n8588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.counter_926__i0_LC_9_14_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i0_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i0_LC_9_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i0_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__31497),
            .in2(_gnd_net_),
            .in3(N__27566),
            .lcout(\Inst_core.Inst_sampler.counter_0 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\Inst_core.Inst_sampler.n7948 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i1_LC_9_14_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i1_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i1_LC_9_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i1_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__30557),
            .in2(_gnd_net_),
            .in3(N__27563),
            .lcout(\Inst_core.Inst_sampler.counter_1 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7948 ),
            .carryout(\Inst_core.Inst_sampler.n7949 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i2_LC_9_14_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i2_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i2_LC_9_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i2_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__30703),
            .in2(_gnd_net_),
            .in3(N__27560),
            .lcout(\Inst_core.Inst_sampler.counter_2 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7949 ),
            .carryout(\Inst_core.Inst_sampler.n7950 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i3_LC_9_14_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i3_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i3_LC_9_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i3_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__30503),
            .in2(_gnd_net_),
            .in3(N__27557),
            .lcout(\Inst_core.Inst_sampler.counter_3 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7950 ),
            .carryout(\Inst_core.Inst_sampler.n7951 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i4_LC_9_14_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i4_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i4_LC_9_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i4_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__27554),
            .in2(_gnd_net_),
            .in3(N__27536),
            .lcout(\Inst_core.Inst_sampler.counter_4 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7951 ),
            .carryout(\Inst_core.Inst_sampler.n7952 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i5_LC_9_14_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i5_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i5_LC_9_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i5_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__32019),
            .in2(_gnd_net_),
            .in3(N__27533),
            .lcout(\Inst_core.Inst_sampler.counter_5 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7952 ),
            .carryout(\Inst_core.Inst_sampler.n7953 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i6_LC_9_14_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i6_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i6_LC_9_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i6_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__31654),
            .in2(_gnd_net_),
            .in3(N__27530),
            .lcout(\Inst_core.Inst_sampler.counter_6 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7953 ),
            .carryout(\Inst_core.Inst_sampler.n7954 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i7_LC_9_14_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i7_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i7_LC_9_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i7_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__27527),
            .in2(_gnd_net_),
            .in3(N__27509),
            .lcout(\Inst_core.Inst_sampler.counter_7 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7954 ),
            .carryout(\Inst_core.Inst_sampler.n7955 ),
            .clk(N__37608),
            .ce(),
            .sr(N__27756));
    defparam \Inst_core.Inst_sampler.counter_926__i8_LC_9_15_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i8_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i8_LC_9_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i8_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__27501),
            .in2(_gnd_net_),
            .in3(N__27479),
            .lcout(\Inst_core.Inst_sampler.counter_8 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\Inst_core.Inst_sampler.n7956 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i9_LC_9_15_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i9_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i9_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i9_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__27700),
            .in2(_gnd_net_),
            .in3(N__27680),
            .lcout(\Inst_core.Inst_sampler.counter_9 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7956 ),
            .carryout(\Inst_core.Inst_sampler.n7957 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i10_LC_9_15_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i10_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i10_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i10_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__27675),
            .in2(_gnd_net_),
            .in3(N__27659),
            .lcout(\Inst_core.Inst_sampler.counter_10 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7957 ),
            .carryout(\Inst_core.Inst_sampler.n7958 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i11_LC_9_15_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i11_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i11_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i11_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__30721),
            .in2(_gnd_net_),
            .in3(N__27656),
            .lcout(\Inst_core.Inst_sampler.counter_11 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7958 ),
            .carryout(\Inst_core.Inst_sampler.n7959 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i12_LC_9_15_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i12_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i12_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i12_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__31549),
            .in2(_gnd_net_),
            .in3(N__27653),
            .lcout(\Inst_core.Inst_sampler.counter_12 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7959 ),
            .carryout(\Inst_core.Inst_sampler.n7960 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i13_LC_9_15_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i13_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i13_LC_9_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i13_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__27650),
            .in2(_gnd_net_),
            .in3(N__27635),
            .lcout(\Inst_core.Inst_sampler.counter_13 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7960 ),
            .carryout(\Inst_core.Inst_sampler.n7961 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i14_LC_9_15_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i14_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i14_LC_9_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i14_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__27632),
            .in2(_gnd_net_),
            .in3(N__27617),
            .lcout(\Inst_core.Inst_sampler.counter_14 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7961 ),
            .carryout(\Inst_core.Inst_sampler.n7962 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i15_LC_9_15_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i15_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i15_LC_9_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i15_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__27614),
            .in2(_gnd_net_),
            .in3(N__27599),
            .lcout(\Inst_core.Inst_sampler.counter_15 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7962 ),
            .carryout(\Inst_core.Inst_sampler.n7963 ),
            .clk(N__37615),
            .ce(),
            .sr(N__27763));
    defparam \Inst_core.Inst_sampler.counter_926__i16_LC_9_16_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i16_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i16_LC_9_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i16_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__27591),
            .in2(_gnd_net_),
            .in3(N__27569),
            .lcout(\Inst_core.Inst_sampler.counter_16 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\Inst_core.Inst_sampler.n7964 ),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_sampler.counter_926__i17_LC_9_16_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i17_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i17_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i17_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__27880),
            .in2(_gnd_net_),
            .in3(N__27860),
            .lcout(\Inst_core.Inst_sampler.counter_17 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7964 ),
            .carryout(\Inst_core.Inst_sampler.n7965 ),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_sampler.counter_926__i18_LC_9_16_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i18_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i18_LC_9_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i18_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__30609),
            .in2(_gnd_net_),
            .in3(N__27857),
            .lcout(\Inst_core.Inst_sampler.counter_18 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7965 ),
            .carryout(\Inst_core.Inst_sampler.n7966 ),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_sampler.counter_926__i19_LC_9_16_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i19_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i19_LC_9_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i19_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__27849),
            .in2(_gnd_net_),
            .in3(N__27827),
            .lcout(\Inst_core.Inst_sampler.counter_19 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7966 ),
            .carryout(\Inst_core.Inst_sampler.n7967 ),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_sampler.counter_926__i20_LC_9_16_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i20_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i20_LC_9_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i20_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__27824),
            .in2(_gnd_net_),
            .in3(N__27809),
            .lcout(\Inst_core.Inst_sampler.counter_20 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7967 ),
            .carryout(\Inst_core.Inst_sampler.n7968 ),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_sampler.counter_926__i21_LC_9_16_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i21_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i21_LC_9_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i21_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__27798),
            .in2(_gnd_net_),
            .in3(N__27776),
            .lcout(\Inst_core.Inst_sampler.counter_21 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7968 ),
            .carryout(\Inst_core.Inst_sampler.n7969 ),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_sampler.counter_926__i22_LC_9_16_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_sampler.counter_926__i22_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i22_LC_9_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i22_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__32080),
            .in2(_gnd_net_),
            .in3(N__27773),
            .lcout(\Inst_core.Inst_sampler.counter_22 ),
            .ltout(),
            .carryin(\Inst_core.Inst_sampler.n7969 ),
            .carryout(\Inst_core.Inst_sampler.n7970 ),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_sampler.counter_926__i23_LC_9_16_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.counter_926__i23_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.counter_926__i23_LC_9_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_sampler.counter_926__i23_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__30745),
            .in2(_gnd_net_),
            .in3(N__27770),
            .lcout(\Inst_core.Inst_sampler.counter_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37622),
            .ce(),
            .sr(N__27767));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.match_84_LC_11_1_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.match_84_LC_11_1_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.match_84_LC_11_1_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.match_84_LC_11_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27728),
            .lcout(\Inst_core.Inst_trigger.stageMatch_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37624),
            .ce(N__32632),
            .sr(N__27710));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.run_83_LC_11_2_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.run_83_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.run_83_LC_11_2_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.run_83_LC_11_2_0  (
            .in0(N__32631),
            .in1(N__32489),
            .in2(N__31862),
            .in3(N__28351),
            .lcout(\Inst_core.stageRun_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37618),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i25_LC_11_2_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i25_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i25_LC_11_2_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i25_LC_11_2_1  (
            .in0(N__28191),
            .in1(_gnd_net_),
            .in2(N__29324),
            .in3(N__31857),
            .lcout(\Inst_core.configRegister_27_adj_1196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37618),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i25_LC_11_2_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i25_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i25_LC_11_2_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i25_LC_11_2_3  (
            .in0(N__28190),
            .in1(N__34105),
            .in2(_gnd_net_),
            .in3(N__32661),
            .lcout(\Inst_core.Inst_trigger.configRegister_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37618),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i1_LC_11_2_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i1_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i1_LC_11_2_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i1_LC_11_2_5  (
            .in0(N__29294),
            .in1(N__35998),
            .in2(_gnd_net_),
            .in3(N__28309),
            .lcout(configRegister_0_adj_1320),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37618),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i1_LC_11_2_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i1_LC_11_2_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i1_LC_11_2_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i1_LC_11_2_6  (
            .in0(N__35999),
            .in1(N__35833),
            .in2(_gnd_net_),
            .in3(N__28132),
            .lcout(configRegister_0_adj_1360),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37618),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i2_LC_11_2_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i2_LC_11_2_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i2_LC_11_2_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i2_LC_11_2_7  (
            .in0(N__29295),
            .in1(N__34268),
            .in2(_gnd_net_),
            .in3(N__28270),
            .lcout(configRegister_1_adj_1319),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37618),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i4_LC_11_3_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i4_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i4_LC_11_3_0 .LUT_INIT=16'b0010011111011000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i4_LC_11_3_0  (
            .in0(N__33556),
            .in1(N__28121),
            .in2(N__28097),
            .in3(N__28865),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37611),
            .ce(),
            .sr(N__27986));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_adj_77_LC_11_3_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_adj_77_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_adj_77_LC_11_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_adj_77_LC_11_3_1  (
            .in0(N__27968),
            .in1(N__27956),
            .in2(N__27947),
            .in3(N__27932),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i5511_2_lut_LC_11_3_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i5511_2_lut_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i5511_2_lut_LC_11_3_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i5511_2_lut_LC_11_3_2  (
            .in0(N__32948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36563),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n6675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_4_lut_LC_11_3_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_4_lut_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_4_lut_LC_11_3_3 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i1_4_lut_LC_11_3_3  (
            .in0(N__36844),
            .in1(N__28339),
            .in2(N__27914),
            .in3(N__27910),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i12_4_lut_LC_11_3_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i12_4_lut_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i12_4_lut_LC_11_3_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i12_4_lut_LC_11_3_4  (
            .in0(N__28789),
            .in1(N__28451),
            .in2(N__28679),
            .in3(N__28394),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7651_2_lut_4_lut_LC_11_3_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7651_2_lut_4_lut_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7651_2_lut_4_lut_LC_11_3_5 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i7651_2_lut_4_lut_LC_11_3_5  (
            .in0(N__36564),
            .in1(N__28338),
            .in2(N__36867),
            .in3(N__32950),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n8626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7561_2_lut_3_lut_LC_11_3_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7561_2_lut_3_lut_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i7561_2_lut_3_lut_LC_11_3_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i7561_2_lut_3_lut_LC_11_3_6  (
            .in0(N__32949),
            .in1(N__36565),
            .in2(_gnd_net_),
            .in3(N__28340),
            .lcout(\Inst_core.n8837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i834_2_lut_3_lut_LC_11_3_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i834_2_lut_3_lut_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i834_2_lut_3_lut_LC_11_3_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i834_2_lut_3_lut_LC_11_3_7  (
            .in0(N__36562),
            .in1(N__28337),
            .in2(_gnd_net_),
            .in3(N__32947),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n1662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i0_LC_11_4_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i0_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i0_LC_11_4_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i0_LC_11_4_0  (
            .in0(N__28310),
            .in1(N__28295),
            .in2(N__33014),
            .in3(N__28280),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_0 ),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7884 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i1_LC_11_4_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i1_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i1_LC_11_4_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i1_LC_11_4_1  (
            .in0(N__28277),
            .in1(N__28710),
            .in2(N__32981),
            .in3(N__28259),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_1 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7884 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7885 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i2_LC_11_4_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i2_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i2_LC_11_4_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i2_LC_11_4_2  (
            .in0(N__28256),
            .in1(N__32912),
            .in2(N__28743),
            .in3(N__28241),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_2 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7885 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7886 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i3_LC_11_4_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i3_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i3_LC_11_4_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i3_LC_11_4_3  (
            .in0(N__28238),
            .in1(N__28714),
            .in2(N__32858),
            .in3(N__28223),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_3 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7886 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7887 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i4_LC_11_4_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i4_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i4_LC_11_4_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i4_LC_11_4_4  (
            .in0(N__28220),
            .in1(N__32995),
            .in2(N__28744),
            .in3(N__28202),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_4 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7887 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7888 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i5_LC_11_4_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i5_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i5_LC_11_4_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i5_LC_11_4_5  (
            .in0(N__28553),
            .in1(N__28718),
            .in2(N__32831),
            .in3(N__28538),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_5 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7888 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7889 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i6_LC_11_4_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i6_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i6_LC_11_4_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i6_LC_11_4_6  (
            .in0(N__28535),
            .in1(N__32240),
            .in2(N__28745),
            .in3(N__28520),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_6 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7889 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7890 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i7_LC_11_4_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i7_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i7_LC_11_4_7 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i7_LC_11_4_7  (
            .in0(N__28517),
            .in1(N__28722),
            .in2(N__32897),
            .in3(N__28496),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_7 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7890 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7891 ),
            .clk(N__37602),
            .ce(N__28657),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i8_LC_11_5_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i8_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i8_LC_11_5_0 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i8_LC_11_5_0  (
            .in0(N__28493),
            .in1(N__28749),
            .in2(N__32813),
            .in3(N__28472),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_8 ),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7892 ),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i9_LC_11_5_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i9_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i9_LC_11_5_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i9_LC_11_5_1  (
            .in0(N__28469),
            .in1(N__28450),
            .in2(N__28766),
            .in3(N__28436),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_9 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7892 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7893 ),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i10_LC_11_5_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i10_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i10_LC_11_5_2 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i10_LC_11_5_2  (
            .in0(N__28433),
            .in1(N__28753),
            .in2(N__32879),
            .in3(N__28415),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_10 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7893 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7894 ),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i11_LC_11_5_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i11_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i11_LC_11_5_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i11_LC_11_5_3  (
            .in0(N__28412),
            .in1(N__28393),
            .in2(N__28767),
            .in3(N__28379),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_11 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7894 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7895 ),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i12_LC_11_5_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i12_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i12_LC_11_5_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i12_LC_11_5_4  (
            .in0(N__28376),
            .in1(N__28757),
            .in2(N__32930),
            .in3(N__28361),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_12 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7895 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7896 ),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i13_LC_11_5_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i13_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i13_LC_11_5_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i13_LC_11_5_5  (
            .in0(N__28811),
            .in1(N__32843),
            .in2(N__28768),
            .in3(N__28793),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_13 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7896 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7897 ),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i14_LC_11_5_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i14_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i14_LC_11_5_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i14_LC_11_5_6  (
            .in0(N__29147),
            .in1(N__28761),
            .in2(N__28790),
            .in3(N__28772),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_14 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7897 ),
            .carryout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n7898 ),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i15_LC_11_5_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i15_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i15_LC_11_5_7 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.counter__i15_LC_11_5_7  (
            .in0(N__28762),
            .in1(N__28675),
            .in2(N__28850),
            .in3(N__28682),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37591),
            .ce(N__28661),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i2_LC_11_6_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i2_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i2_LC_11_6_0 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i2_LC_11_6_0  (
            .in0(N__28646),
            .in1(N__33552),
            .in2(N__29573),
            .in3(N__30928),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37578),
            .ce(),
            .sr(N__28622));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i11_4_lut_LC_11_6_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i11_4_lut_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i11_4_lut_LC_11_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i11_4_lut_LC_11_6_1  (
            .in0(N__33859),
            .in1(N__32737),
            .in2(N__33151),
            .in3(N__33061),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i12_4_lut_LC_11_6_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i12_4_lut_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i12_4_lut_LC_11_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i12_4_lut_LC_11_6_2  (
            .in0(N__33799),
            .in1(N__33097),
            .in2(N__33709),
            .in3(N__33028),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_2_lut_LC_11_6_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_2_lut_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_2_lut_LC_11_6_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_2_lut_LC_11_6_3  (
            .in0(N__35084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28963),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i44_4_lut_LC_11_6_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i44_4_lut_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i44_4_lut_LC_11_6_4 .LUT_INIT=16'b0100110100000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i44_4_lut_LC_11_6_4  (
            .in0(N__29414),
            .in1(N__28913),
            .in2(N__28607),
            .in3(N__28604),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n100 ),
            .ltout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i133_2_lut_LC_11_6_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i133_2_lut_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i133_2_lut_LC_11_6_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i133_2_lut_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28577),
            .in3(N__28574),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.LessThan_42_i4_4_lut_LC_11_6_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.LessThan_42_i4_4_lut_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.LessThan_42_i4_4_lut_LC_11_6_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.LessThan_42_i4_4_lut_LC_11_6_6  (
            .in0(N__28964),
            .in1(N__28928),
            .in2(N__36125),
            .in3(N__28912),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i4_LC_11_7_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i4_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i4_LC_11_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i4_LC_11_7_0  (
            .in0(N__29130),
            .in1(N__28861),
            .in2(_gnd_net_),
            .in3(N__36092),
            .lcout(valueRegister_4_adj_1372),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i6_LC_11_7_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i6_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i6_LC_11_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i6_LC_11_7_1  (
            .in0(N__34100),
            .in1(N__33202),
            .in2(_gnd_net_),
            .in3(N__31322),
            .lcout(configRegister_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i12_LC_11_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i12_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i12_LC_11_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i12_LC_11_7_2  (
            .in0(N__35310),
            .in1(N__31091),
            .in2(_gnd_net_),
            .in3(N__31524),
            .lcout(divider_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i1_LC_11_7_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i1_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i1_LC_11_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i1_LC_11_7_3  (
            .in0(N__34099),
            .in1(N__35957),
            .in2(_gnd_net_),
            .in3(N__32788),
            .lcout(configRegister_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i16_LC_11_7_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i16_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i16_LC_11_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i16_LC_11_7_4  (
            .in0(N__29292),
            .in1(N__33936),
            .in2(_gnd_net_),
            .in3(N__28843),
            .lcout(configRegister_15_adj_1305),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i7_LC_11_7_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i7_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i7_LC_11_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i7_LC_11_7_5  (
            .in0(N__34101),
            .in1(N__33184),
            .in2(_gnd_net_),
            .in3(N__34421),
            .lcout(configRegister_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i15_LC_11_7_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i15_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i15_LC_11_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i15_LC_11_7_6  (
            .in0(N__35432),
            .in1(N__33935),
            .in2(_gnd_net_),
            .in3(N__28825),
            .lcout(bwd_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i24_LC_11_7_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i24_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i24_LC_11_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i24_LC_11_7_7  (
            .in0(N__29293),
            .in1(N__30296),
            .in2(_gnd_net_),
            .in3(N__35676),
            .lcout(configRegister_26_adj_1297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i18_LC_11_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i18_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i18_LC_11_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i18_LC_11_8_0  (
            .in0(N__29528),
            .in1(N__34104),
            .in2(_gnd_net_),
            .in3(N__29413),
            .lcout(configRegister_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i13_LC_11_8_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i13_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i13_LC_11_8_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i13_LC_11_8_1  (
            .in0(N__29395),
            .in1(N__35433),
            .in2(_gnd_net_),
            .in3(N__29914),
            .lcout(bwd_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i2_LC_11_8_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i2_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i2_LC_11_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i2_LC_11_8_2  (
            .in0(N__34528),
            .in1(N__29692),
            .in2(_gnd_net_),
            .in3(N__29824),
            .lcout(valueRegister_2_adj_1294),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i12_LC_11_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i12_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i12_LC_11_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i12_LC_11_8_3  (
            .in0(N__34102),
            .in1(N__34569),
            .in2(_gnd_net_),
            .in3(N__33040),
            .lcout(configRegister_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i15_LC_11_8_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i15_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i15_LC_11_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.configRegister__i15_LC_11_8_4  (
            .in0(N__29143),
            .in1(N__29291),
            .in2(_gnd_net_),
            .in3(N__30085),
            .lcout(configRegister_14_adj_1306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i5_LC_11_8_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i5_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i5_LC_11_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i5_LC_11_8_5  (
            .in0(N__34103),
            .in1(N__33220),
            .in2(_gnd_net_),
            .in3(N__29131),
            .lcout(configRegister_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i6_LC_11_8_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i6_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i6_LC_11_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i6_LC_11_8_6  (
            .in0(N__34430),
            .in1(N__31092),
            .in2(_gnd_net_),
            .in3(N__30522),
            .lcout(divider_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i1_LC_11_8_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i1_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i1_LC_11_8_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i1_LC_11_8_7  (
            .in0(N__36099),
            .in1(N__34259),
            .in2(_gnd_net_),
            .in3(N__33664),
            .lcout(valueRegister_1_adj_1375),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i14_LC_11_9_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i14_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i14_LC_11_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i14_LC_11_9_0  (
            .in0(N__35506),
            .in1(N__30069),
            .in2(_gnd_net_),
            .in3(N__29848),
            .lcout(\Inst_core.Inst_controller.bwd_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i7_LC_11_9_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i7_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i7_LC_11_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i7_LC_11_9_1  (
            .in0(N__35507),
            .in1(N__29764),
            .in2(_gnd_net_),
            .in3(N__28978),
            .lcout(fwd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i1_LC_11_9_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i1_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i1_LC_11_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i1_LC_11_9_2  (
            .in0(N__34262),
            .in1(N__31090),
            .in2(_gnd_net_),
            .in3(N__30636),
            .lcout(divider_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i6_LC_11_9_3 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i6_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i6_LC_11_9_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i6_LC_11_9_3  (
            .in0(N__34431),
            .in1(N__34825),
            .in2(N__31324),
            .in3(N__35052),
            .lcout(cmd_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3592_1_lut_LC_11_9_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3592_1_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i3592_1_lut_LC_11_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i3592_1_lut_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29780),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n4751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i23_LC_11_9_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i23_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i23_LC_11_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i23_LC_11_9_5  (
            .in0(N__31089),
            .in1(N__29765),
            .in2(_gnd_net_),
            .in3(N__30666),
            .lcout(divider_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i2_LC_11_9_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i2_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i2_LC_11_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i2_LC_11_9_7  (
            .in0(N__36090),
            .in1(N__29671),
            .in2(_gnd_net_),
            .in3(N__29566),
            .lcout(valueRegister_2_adj_1374),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i19_LC_11_10_0 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i19_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i19_LC_11_10_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i19_LC_11_10_0  (
            .in0(N__35048),
            .in1(N__30001),
            .in2(N__30034),
            .in3(N__34846),
            .lcout(cmd_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i18_LC_11_10_1 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i18_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i18_LC_11_10_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i18_LC_11_10_1  (
            .in0(N__34843),
            .in1(N__29513),
            .in2(N__30033),
            .in3(N__35049),
            .lcout(cmd_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i17_LC_11_10_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i17_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i17_LC_11_10_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i17_LC_11_10_2  (
            .in0(N__35047),
            .in1(N__36146),
            .in2(N__29527),
            .in3(N__34845),
            .lcout(cmd_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i0_LC_11_10_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i0_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i0_LC_11_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.valueRegister_i0_i0_LC_11_10_3  (
            .in0(N__29489),
            .in1(N__35989),
            .in2(_gnd_net_),
            .in3(N__32209),
            .lcout(valueRegister_0_adj_1336),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i15_LC_11_10_4 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i15_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i15_LC_11_10_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i15_LC_11_10_4  (
            .in0(N__35046),
            .in1(N__30068),
            .in2(N__33941),
            .in3(N__34844),
            .lcout(cmd_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.fwd_i0_i2_LC_11_10_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.fwd_i0_i2_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.fwd_i0_i2_LC_11_10_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_controller.fwd_i0_i2_LC_11_10_5  (
            .in0(N__30023),
            .in1(N__35508),
            .in2(_gnd_net_),
            .in3(N__30187),
            .lcout(fwd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i19_LC_11_10_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i19_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i19_LC_11_10_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i19_LC_11_10_7  (
            .in0(N__31093),
            .in1(_gnd_net_),
            .in2(N__30002),
            .in3(N__29958),
            .lcout(divider_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_62_LC_11_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_62_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1_4_lut_adj_62_LC_11_11_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \Inst_core.Inst_controller.i1_4_lut_adj_62_LC_11_11_0  (
            .in0(N__37723),
            .in1(N__29936),
            .in2(N__29918),
            .in3(N__37099),
            .lcout(),
            .ltout(\Inst_core.Inst_controller.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i13_4_lut_LC_11_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i13_4_lut_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i13_4_lut_LC_11_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_controller.i13_4_lut_LC_11_11_1  (
            .in0(N__29900),
            .in1(N__29888),
            .in2(N__29879),
            .in3(N__29834),
            .lcout(),
            .ltout(\Inst_core.Inst_controller.n29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i1_3_lut_4_lut_LC_11_11_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1_3_lut_4_lut_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1_3_lut_4_lut_LC_11_11_2 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \Inst_core.Inst_controller.i1_3_lut_4_lut_LC_11_11_2  (
            .in0(N__36274),
            .in1(N__29876),
            .in2(N__29864),
            .in3(N__36256),
            .lcout(\Inst_core.Inst_controller.nstate_1_N_827_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i5529_2_lut_LC_11_11_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i5529_2_lut_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i5529_2_lut_LC_11_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_core.Inst_controller.i5529_2_lut_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__36255),
            .in2(_gnd_net_),
            .in3(N__36273),
            .lcout(\Inst_core.Inst_controller.n6693 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i3_4_lut_adj_61_LC_11_11_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i3_4_lut_adj_61_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i3_4_lut_adj_61_LC_11_11_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_controller.i3_4_lut_adj_61_LC_11_11_4  (
            .in0(N__29849),
            .in1(N__37696),
            .in2(N__35873),
            .in3(N__36235),
            .lcout(\Inst_core.Inst_controller.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i2_LC_11_11_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i2_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i2_LC_11_11_5 .LUT_INIT=16'b0110011001011010;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i2_LC_11_11_5  (
            .in0(N__29828),
            .in1(N__29813),
            .in2(N__30941),
            .in3(N__30344),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37590),
            .ce(),
            .sr(N__30482));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i6_LC_11_12_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i6_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i6_LC_11_12_0 .LUT_INIT=16'b0011011011000110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_i6_LC_11_12_0  (
            .in0(N__30442),
            .in1(N__34301),
            .in2(N__30347),
            .in3(N__30254),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.intermediateRegister_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37601),
            .ce(),
            .sr(N__30221));
    defparam \Inst_core.Inst_controller.i4_4_lut_LC_11_12_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i4_4_lut_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i4_4_lut_LC_11_12_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_controller.i4_4_lut_LC_11_12_1  (
            .in0(N__30209),
            .in1(N__37098),
            .in2(N__30191),
            .in3(N__36234),
            .lcout(\Inst_core.Inst_controller.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i102_2_lut_LC_11_12_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i102_2_lut_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i102_2_lut_LC_11_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_core.Inst_controller.i102_2_lut_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__36447),
            .in2(_gnd_net_),
            .in3(N__36317),
            .lcout(debugleds_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_decoder.i1_2_lut_LC_11_12_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_decoder.i1_2_lut_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_decoder.i1_2_lut_LC_11_12_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Inst_core.Inst_decoder.i1_2_lut_LC_11_12_3  (
            .in0(N__36448),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36871),
            .lcout(),
            .ltout(\Inst_core.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i7628_4_lut_LC_11_12_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i7628_4_lut_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i7628_4_lut_LC_11_12_4 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \Inst_core.Inst_controller.i7628_4_lut_LC_11_12_4  (
            .in0(N__36512),
            .in1(N__30144),
            .in2(N__30125),
            .in3(N__36674),
            .lcout(\Inst_core.Inst_controller.n3907 ),
            .ltout(\Inst_core.Inst_controller.n3907_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i7641_4_lut_LC_11_12_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i7641_4_lut_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i7641_4_lut_LC_11_12_5 .LUT_INIT=16'b0010000011110000;
    LogicCell40 \Inst_core.Inst_controller.i7641_4_lut_LC_11_12_5  (
            .in0(N__36318),
            .in1(N__35184),
            .in2(N__30122),
            .in3(N__36281),
            .lcout(\Inst_core.Inst_controller.n4691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i7666_3_lut_4_lut_LC_11_12_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i7666_3_lut_4_lut_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i7666_3_lut_4_lut_LC_11_12_6 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i7666_3_lut_4_lut_LC_11_12_6  (
            .in0(N__33267),
            .in1(N__32450),
            .in2(N__36553),
            .in3(N__36872),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7668_1_lut_2_lut_3_lut_LC_11_12_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7668_1_lut_2_lut_3_lut_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7668_1_lut_2_lut_3_lut_LC_11_12_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Inst_core.Inst_sampler.i7668_1_lut_2_lut_3_lut_LC_11_12_7  (
            .in0(N__32449),
            .in1(N__36508),
            .in2(_gnd_net_),
            .in3(N__33266),
            .lcout(\Inst_core.n9053 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i2_LC_11_13_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i2_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i2_LC_11_13_0 .LUT_INIT=16'b0011011011000110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i2_LC_11_13_0  (
            .in0(N__30940),
            .in1(N__30845),
            .in2(N__35578),
            .in3(N__30827),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37610),
            .ce(),
            .sr(N__30803));
    defparam \Inst_core.Inst_sampler.i12_4_lut_LC_11_13_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i12_4_lut_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i12_4_lut_LC_11_13_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_sampler.i12_4_lut_LC_11_13_1  (
            .in0(N__30784),
            .in1(N__30727),
            .in2(N__30671),
            .in3(N__30749),
            .lcout(\Inst_core.Inst_sampler.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7250_4_lut_LC_11_13_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7250_4_lut_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7250_4_lut_LC_11_13_2 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \Inst_core.Inst_sampler.i7250_4_lut_LC_11_13_2  (
            .in0(N__31505),
            .in1(N__30638),
            .in2(N__30731),
            .in3(N__31528),
            .lcout(\Inst_core.Inst_sampler.n8618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.counter_22__I_0_i3_2_lut_LC_11_13_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.counter_22__I_0_i3_2_lut_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.counter_22__I_0_i3_2_lut_LC_11_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Inst_core.Inst_sampler.counter_22__I_0_i3_2_lut_LC_11_13_3  (
            .in0(N__31687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30707),
            .lcout(),
            .ltout(\Inst_core.Inst_sampler.n3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7288_4_lut_LC_11_13_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7288_4_lut_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7288_4_lut_LC_11_13_4 .LUT_INIT=16'b1111101111111110;
    LogicCell40 \Inst_core.Inst_sampler.i7288_4_lut_LC_11_13_4  (
            .in0(N__30683),
            .in1(N__30524),
            .in2(N__30674),
            .in3(N__32027),
            .lcout(),
            .ltout(\Inst_core.Inst_sampler.n8656_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7304_4_lut_LC_11_13_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7304_4_lut_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7304_4_lut_LC_11_13_5 .LUT_INIT=16'b1111110111111110;
    LogicCell40 \Inst_core.Inst_sampler.i7304_4_lut_LC_11_13_5  (
            .in0(N__30670),
            .in1(N__30650),
            .in2(N__30641),
            .in3(N__32081),
            .lcout(\Inst_core.Inst_sampler.n8673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i3_4_lut_LC_11_14_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i3_4_lut_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i3_4_lut_LC_11_14_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i3_4_lut_LC_11_14_0  (
            .in0(N__30637),
            .in1(N__30616),
            .in2(N__30590),
            .in3(N__30556),
            .lcout(),
            .ltout(\Inst_core.Inst_sampler.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i19_4_lut_LC_11_14_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i19_4_lut_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i19_4_lut_LC_11_14_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_sampler.i19_4_lut_LC_11_14_1  (
            .in0(N__30536),
            .in1(N__31631),
            .in2(N__30527),
            .in3(N__31478),
            .lcout(\Inst_core.Inst_sampler.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i2_4_lut_LC_11_14_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i2_4_lut_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i2_4_lut_LC_11_14_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i2_4_lut_LC_11_14_2  (
            .in0(N__30523),
            .in1(N__30502),
            .in2(N__31688),
            .in3(N__31650),
            .lcout(\Inst_core.Inst_sampler.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i3_LC_11_14_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i3_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i3_LC_11_14_3 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i3_LC_11_14_3  (
            .in0(N__31625),
            .in1(N__31604),
            .in2(N__35610),
            .in3(N__32352),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37617),
            .ce(),
            .sr(N__31583));
    defparam \Inst_core.Inst_sampler.i1_4_lut_LC_11_14_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i1_4_lut_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i1_4_lut_LC_11_14_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i1_4_lut_LC_11_14_4  (
            .in0(N__31568),
            .in1(N__31553),
            .in2(N__31529),
            .in3(N__31498),
            .lcout(\Inst_core.Inst_sampler.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i7_LC_11_15_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i7_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.Inst_filter.input360_i7_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Inst_core.Inst_sync.Inst_filter.input360_i7_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31428),
            .lcout(\Inst_core.Inst_sync.Inst_filter.input360_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37623),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sync.synchronizedInput_i7_LC_11_15_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_sync.synchronizedInput_i7_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sync.synchronizedInput_i7_LC_11_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Inst_core.Inst_sync.synchronizedInput_i7_LC_11_15_1  (
            .in0(N__31460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Inst_core.Inst_sync.synchronizedInput_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37623),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.divider_i0_i5_LC_11_15_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.divider_i0_i5_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.divider_i0_i5_LC_11_15_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_sampler.divider_i0_i5_LC_11_15_2  (
            .in0(N__31323),
            .in1(N__31103),
            .in2(_gnd_net_),
            .in3(N__32101),
            .lcout(divider_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37623),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i21_4_lut_LC_11_15_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i21_4_lut_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i21_4_lut_LC_11_15_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_sampler.i21_4_lut_LC_11_15_3  (
            .in0(N__31997),
            .in1(N__31232),
            .in2(N__31223),
            .in3(N__31211),
            .lcout(\Inst_core.Inst_sampler.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.ready_40_LC_11_15_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.ready_40_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_sampler.ready_40_LC_11_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Inst_core.Inst_sampler.ready_40_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__31102),
            .in2(_gnd_net_),
            .in3(N__31896),
            .lcout(sampleReady),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37623),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7611_4_lut_LC_11_15_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7611_4_lut_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7611_4_lut_LC_11_15_5 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \Inst_core.Inst_sampler.i7611_4_lut_LC_11_15_5  (
            .in0(N__31895),
            .in1(N__30974),
            .in2(N__30962),
            .in3(N__30950),
            .lcout(\Inst_core.Inst_sampler.n8687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i0_LC_11_16_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i0_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i0_LC_11_16_0 .LUT_INIT=16'b0110010101101010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_i0_LC_11_16_0  (
            .in0(N__32213),
            .in1(N__32198),
            .in2(N__35605),
            .in3(N__31800),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.intermediateRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37627),
            .ce(),
            .sr(N__32177));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_LC_11_16_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_LC_11_16_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.i3_4_lut_LC_11_16_1  (
            .in0(N__32162),
            .in1(N__32150),
            .in2(N__32141),
            .in3(N__32129),
            .lcout(\Inst_core.Inst_trigger.stages_2__Inst_stage.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i10_4_lut_LC_11_16_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i10_4_lut_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i10_4_lut_LC_11_16_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \Inst_core.Inst_sampler.i10_4_lut_LC_11_16_2  (
            .in0(N__32097),
            .in1(N__32076),
            .in2(N__32057),
            .in3(N__32026),
            .lcout(\Inst_core.Inst_sampler.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i7609_3_lut_LC_11_16_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i7609_3_lut_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i7609_3_lut_LC_11_16_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Inst_core.Inst_sampler.i7609_3_lut_LC_11_16_4  (
            .in0(N__31991),
            .in1(N__31979),
            .in2(_gnd_net_),
            .in3(N__31970),
            .lcout(ready50_N_581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.match_84_LC_12_1_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.match_84_LC_12_1_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.match_84_LC_12_1_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.match_84_LC_12_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31861),
            .lcout(\Inst_core.Inst_trigger.stageMatch_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37628),
            .ce(N__32620),
            .sr(N__31844));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.match_84_LC_12_2_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.match_84_LC_12_2_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.match_84_LC_12_2_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.match_84_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32662),
            .lcout(\Inst_core.Inst_trigger.stageMatch_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37626),
            .ce(N__32639),
            .sr(N__31832));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i0_LC_12_3_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i0_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i0_LC_12_3_0 .LUT_INIT=16'b0101011010011010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i0_LC_12_3_0  (
            .in0(N__36020),
            .in1(N__33559),
            .in2(N__31804),
            .in3(N__31715),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37620),
            .ce(),
            .sr(N__32705));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_LC_12_3_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_LC_12_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i3_4_lut_LC_12_3_1  (
            .in0(N__33443),
            .in1(N__32693),
            .in2(N__32264),
            .in3(N__32681),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7_adj_1000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_76_LC_12_3_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_76_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_76_LC_12_3_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i1_2_lut_adj_76_LC_12_3_2  (
            .in0(N__33259),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36612),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n8521_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i18_4_lut_LC_12_3_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i18_4_lut_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.i18_4_lut_LC_12_3_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.i18_4_lut_LC_12_3_3  (
            .in0(N__32663),
            .in1(N__32542),
            .in2(N__32642),
            .in3(N__32621),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.i3_4_lut_LC_12_3_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.i3_4_lut_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.i3_4_lut_LC_12_3_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.i3_4_lut_LC_12_3_4  (
            .in0(N__32543),
            .in1(N__32528),
            .in2(N__32510),
            .in3(N__32488),
            .lcout(\Inst_core.nstate_1_N_831_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i7508_2_lut_LC_12_3_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i7508_2_lut_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i7508_2_lut_LC_12_3_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i7508_2_lut_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__36611),
            .in2(_gnd_net_),
            .in3(N__33260),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n8753_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_4_lut_LC_12_3_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_4_lut_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_4_lut_LC_12_3_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i1_4_lut_LC_12_3_6  (
            .in0(N__32439),
            .in1(N__36866),
            .in2(N__32477),
            .in3(N__32473),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n4044 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_sampler.i1_2_lut_3_lut_LC_12_3_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_sampler.i1_2_lut_3_lut_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_sampler.i1_2_lut_3_lut_LC_12_3_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Inst_core.Inst_sampler.i1_2_lut_3_lut_LC_12_3_7  (
            .in0(N__32438),
            .in1(N__36610),
            .in2(_gnd_net_),
            .in3(N__33258),
            .lcout(\Inst_core.n1705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i3_LC_12_4_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i3_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i3_LC_12_4_0 .LUT_INIT=16'b0110011001011010;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i3_LC_12_4_0  (
            .in0(N__32396),
            .in1(N__32381),
            .in2(N__32360),
            .in3(N__33558),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37613),
            .ce(),
            .sr(N__32255));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i9_4_lut_LC_12_4_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i9_4_lut_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i9_4_lut_LC_12_4_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i9_4_lut_LC_12_4_1  (
            .in0(N__32239),
            .in1(N__33010),
            .in2(N__32999),
            .in3(N__32977),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i15_4_lut_LC_12_4_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i15_4_lut_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i15_4_lut_LC_12_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i15_4_lut_LC_12_4_2  (
            .in0(N__32966),
            .in1(N__32798),
            .in2(N__32960),
            .in3(N__32864),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i11_4_lut_LC_12_4_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i11_4_lut_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i11_4_lut_LC_12_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i11_4_lut_LC_12_4_3  (
            .in0(N__32929),
            .in1(N__32908),
            .in2(N__32896),
            .in3(N__32875),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i10_4_lut_LC_12_4_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i10_4_lut_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.i10_4_lut_LC_12_4_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.i10_4_lut_LC_12_4_4  (
            .in0(N__32854),
            .in1(N__32842),
            .in2(N__32830),
            .in3(N__32809),
            .lcout(\Inst_core.Inst_trigger.stages_1__Inst_stage.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i0_LC_12_5_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i0_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i0_LC_12_5_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i0_LC_12_5_0  (
            .in0(N__32792),
            .in1(N__32777),
            .in2(N__33302),
            .in3(N__32765),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_0 ),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7869 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i1_LC_12_5_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i1_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i1_LC_12_5_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i1_LC_12_5_1  (
            .in0(N__35099),
            .in1(N__33753),
            .in2(N__33338),
            .in3(N__32762),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_1 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7869 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7870 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i2_LC_12_5_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i2_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i2_LC_12_5_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i2_LC_12_5_2  (
            .in0(N__32759),
            .in1(N__32738),
            .in2(N__33780),
            .in3(N__32726),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_2 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7870 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7871 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i3_LC_12_5_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i3_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i3_LC_12_5_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i3_LC_12_5_3  (
            .in0(N__32723),
            .in1(N__33757),
            .in2(N__35123),
            .in3(N__32708),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_3 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7871 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7872 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i4_LC_12_5_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i4_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i4_LC_12_5_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i4_LC_12_5_4  (
            .in0(N__33224),
            .in1(N__33316),
            .in2(N__33781),
            .in3(N__33209),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_4 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7872 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7873 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i5_LC_12_5_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i5_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i5_LC_12_5_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i5_LC_12_5_5  (
            .in0(N__33206),
            .in1(N__33761),
            .in2(N__35143),
            .in3(N__33191),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_5 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7873 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7874 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i6_LC_12_5_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i6_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i6_LC_12_5_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i6_LC_12_5_6  (
            .in0(N__33188),
            .in1(N__33352),
            .in2(N__33782),
            .in3(N__33173),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_6 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7874 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7875 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i7_LC_12_5_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i7_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i7_LC_12_5_7 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i7_LC_12_5_7  (
            .in0(N__33170),
            .in1(N__33765),
            .in2(N__33152),
            .in3(N__33134),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_7 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7875 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7876 ),
            .clk(N__37604),
            .ce(N__33692),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i8_LC_12_6_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i8_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i8_LC_12_6_0 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i8_LC_12_6_0  (
            .in0(N__33131),
            .in1(N__33766),
            .in2(N__35171),
            .in3(N__33116),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_8 ),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7877 ),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i9_LC_12_6_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i9_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i9_LC_12_6_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i9_LC_12_6_1  (
            .in0(N__33113),
            .in1(N__33098),
            .in2(N__33783),
            .in3(N__33086),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_9 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7877 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7878 ),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i10_LC_12_6_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i10_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i10_LC_12_6_2 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i10_LC_12_6_2  (
            .in0(N__33083),
            .in1(N__33770),
            .in2(N__33065),
            .in3(N__33050),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_10 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7878 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7879 ),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i11_LC_12_6_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i11_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i11_LC_12_6_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i11_LC_12_6_3  (
            .in0(N__33047),
            .in1(N__33029),
            .in2(N__33784),
            .in3(N__33017),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_11 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7879 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7880 ),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i12_LC_12_6_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i12_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i12_LC_12_6_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i12_LC_12_6_4  (
            .in0(N__34283),
            .in1(N__33774),
            .in2(N__33863),
            .in3(N__33848),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_12 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7880 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7881 ),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i13_LC_12_6_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i13_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i13_LC_12_6_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i13_LC_12_6_5  (
            .in0(N__33845),
            .in1(N__35156),
            .in2(N__33785),
            .in3(N__33824),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_13 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7881 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7882 ),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i14_LC_12_6_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i14_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i14_LC_12_6_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i14_LC_12_6_6  (
            .in0(N__33821),
            .in1(N__33778),
            .in2(N__33803),
            .in3(N__33788),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_14 ),
            .ltout(),
            .carryin(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7882 ),
            .carryout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n7883 ),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i15_LC_12_6_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i15_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i15_LC_12_6_7 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.counter__i15_LC_12_6_7  (
            .in0(N__33779),
            .in1(N__33878),
            .in2(N__33710),
            .in3(N__33713),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37593),
            .ce(N__33691),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i1_LC_12_7_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i1_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i1_LC_12_7_0 .LUT_INIT=16'b0101011010100110;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_i1_LC_12_7_0  (
            .in0(N__33668),
            .in1(N__33647),
            .in2(N__33560),
            .in3(N__33467),
            .lcout(\Inst_core.Inst_trigger.stages_3__Inst_stage.intermediateRegister_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37579),
            .ce(),
            .sr(N__33431));
    defparam \Inst_core.Inst_trigger.i3_4_lut_adj_78_LC_12_7_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.i3_4_lut_adj_78_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.i3_4_lut_adj_78_LC_12_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.i3_4_lut_adj_78_LC_12_7_1  (
            .in0(N__33419),
            .in1(N__33404),
            .in2(N__33392),
            .in3(N__33377),
            .lcout(\Inst_core.Inst_trigger.levelReg_1__N_590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i9_4_lut_LC_12_7_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i9_4_lut_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i9_4_lut_LC_12_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i9_4_lut_LC_12_7_2  (
            .in0(N__33353),
            .in1(N__33337),
            .in2(N__33320),
            .in3(N__33301),
            .lcout(),
            .ltout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i15_4_lut_LC_12_7_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i15_4_lut_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i15_4_lut_LC_12_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i15_4_lut_LC_12_7_3  (
            .in0(N__33284),
            .in1(N__35105),
            .in2(N__33278),
            .in3(N__33275),
            .lcout(\Inst_core.n31_adj_1132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i10_4_lut_LC_12_7_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i10_4_lut_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.i10_4_lut_LC_12_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.i10_4_lut_LC_12_7_4  (
            .in0(N__35167),
            .in1(N__35155),
            .in2(N__35144),
            .in3(N__35122),
            .lcout(\Inst_core.Inst_trigger.stages_0__Inst_stage.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i2_LC_12_8_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i2_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i2_LC_12_8_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i2_LC_12_8_0  (
            .in0(N__34261),
            .in1(_gnd_net_),
            .in2(N__34124),
            .in3(N__35095),
            .lcout(configRegister_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i17_LC_12_8_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i17_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i17_LC_12_8_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i17_LC_12_8_1  (
            .in0(N__36160),
            .in1(N__34115),
            .in2(_gnd_net_),
            .in3(N__35083),
            .lcout(configRegister_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_eia232.Inst_receiver.dataBuf_i12_LC_12_8_2 .C_ON=1'b0;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i12_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \Inst_eia232.Inst_receiver.dataBuf_i12_LC_12_8_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \Inst_eia232.Inst_receiver.dataBuf_i12_LC_12_8_2  (
            .in0(N__34568),
            .in1(N__34964),
            .in2(N__34850),
            .in3(N__35312),
            .lcout(cmd_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i6_LC_12_8_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i6_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i6_LC_12_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_1__Inst_stage.valueRegister_i0_i6_LC_12_8_3  (
            .in0(N__34520),
            .in1(N__34432),
            .in2(_gnd_net_),
            .in3(N__34294),
            .lcout(valueRegister_6_adj_1290),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i13_LC_12_8_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i13_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i13_LC_12_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i13_LC_12_8_4  (
            .in0(N__34113),
            .in1(N__35311),
            .in2(_gnd_net_),
            .in3(N__34279),
            .lcout(configRegister_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i1_LC_12_8_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i1_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i1_LC_12_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i1_LC_12_8_5  (
            .in0(N__35505),
            .in1(N__34260),
            .in2(_gnd_net_),
            .in3(N__34138),
            .lcout(bwd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i16_LC_12_8_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i16_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i16_LC_12_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_0__Inst_stage.configRegister__i16_LC_12_8_6  (
            .in0(N__34114),
            .in1(N__33940),
            .in2(_gnd_net_),
            .in3(N__33874),
            .lcout(configRegister_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i17_LC_12_8_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i17_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i17_LC_12_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i17_LC_12_8_7  (
            .in0(N__36161),
            .in1(N__35849),
            .in2(_gnd_net_),
            .in3(N__36118),
            .lcout(configRegister_16_adj_1344),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i0_LC_12_9_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i0_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i0_LC_12_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_trigger.stages_3__Inst_stage.valueRegister_i0_i0_LC_12_9_7  (
            .in0(N__36091),
            .in1(N__35995),
            .in2(_gnd_net_),
            .in3(N__36010),
            .lcout(valueRegister_0_adj_1376),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37580),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i0_LC_12_10_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i0_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i0_LC_12_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i0_LC_12_10_1  (
            .in0(N__35442),
            .in1(N__35996),
            .in2(_gnd_net_),
            .in3(N__35872),
            .lcout(bwd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37592),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i24_LC_12_10_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i24_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i24_LC_12_10_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Inst_core.Inst_trigger.stages_2__Inst_stage.configRegister__i24_LC_12_10_2  (
            .in0(N__35539),
            .in1(N__35848),
            .in2(_gnd_net_),
            .in3(N__35681),
            .lcout(configRegister_26_adj_1337),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37592),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.bwd_i0_i12_LC_12_10_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.bwd_i0_i12_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.bwd_i0_i12_LC_12_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Inst_core.Inst_controller.bwd_i0_i12_LC_12_10_4  (
            .in0(N__35443),
            .in1(N__35309),
            .in2(_gnd_net_),
            .in3(N__35233),
            .lcout(bwd_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37592),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.state_FSM_i2_LC_12_11_0 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.state_FSM_i2_LC_12_11_0 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_controller.state_FSM_i2_LC_12_11_0 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \Inst_core.Inst_controller.state_FSM_i2_LC_12_11_0  (
            .in0(N__36450),
            .in1(N__36705),
            .in2(N__36716),
            .in3(N__36689),
            .lcout(send),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37603),
            .ce(),
            .sr(N__36875));
    defparam \Inst_core.Inst_controller.state_FSM_i1_LC_12_11_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.state_FSM_i1_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_controller.state_FSM_i1_LC_12_11_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Inst_core.Inst_controller.state_FSM_i1_LC_12_11_1  (
            .in0(N__36688),
            .in1(N__35197),
            .in2(N__36707),
            .in3(N__35219),
            .lcout(\Inst_core.Inst_controller.n320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37603),
            .ce(),
            .sr(N__36875));
    defparam \Inst_core.Inst_controller.state_FSM_i0_LC_12_11_2 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.state_FSM_i0_LC_12_11_2 .SEQ_MODE=4'b1011;
    defparam \Inst_core.Inst_controller.state_FSM_i0_LC_12_11_2 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \Inst_core.Inst_controller.state_FSM_i0_LC_12_11_2  (
            .in0(N__36321),
            .in1(N__35215),
            .in2(N__35198),
            .in3(N__35185),
            .lcout(\Inst_core.Inst_controller.n321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37603),
            .ce(),
            .sr(N__36875));
    defparam \Inst_core.Inst_controller.state_FSM_i3_LC_12_11_3 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.state_FSM_i3_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \Inst_core.Inst_controller.state_FSM_i3_LC_12_11_3 .LUT_INIT=16'b1111110010100000;
    LogicCell40 \Inst_core.Inst_controller.state_FSM_i3_LC_12_11_3  (
            .in0(N__35186),
            .in1(N__36731),
            .in2(N__36339),
            .in3(N__36451),
            .lcout(\Inst_core.n318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37603),
            .ce(),
            .sr(N__36875));
    defparam \Inst_core.Inst_controller.i1605_3_lut_LC_12_11_4 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1605_3_lut_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1605_3_lut_LC_12_11_4 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \Inst_core.Inst_controller.i1605_3_lut_LC_12_11_4  (
            .in0(N__36452),
            .in1(N__36325),
            .in2(_gnd_net_),
            .in3(N__36706),
            .lcout(debugleds_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i5479_2_lut_LC_12_11_5 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i5479_2_lut_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i5479_2_lut_LC_12_11_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Inst_core.Inst_controller.i5479_2_lut_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__36730),
            .in2(_gnd_net_),
            .in3(N__36320),
            .lcout(\Inst_core.Inst_controller.nstate_1_N_825_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i1608_2_lut_LC_12_11_6 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i1608_2_lut_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i1608_2_lut_LC_12_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Inst_core.Inst_controller.i1608_2_lut_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__36701),
            .in2(_gnd_net_),
            .in3(N__36687),
            .lcout(\Inst_core.Inst_controller.n2717 ),
            .ltout(\Inst_core.Inst_controller.n2717_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.i5504_3_lut_4_lut_LC_12_11_7 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.i5504_3_lut_4_lut_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \Inst_core.Inst_controller.i5504_3_lut_4_lut_LC_12_11_7 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Inst_core.Inst_controller.i5504_3_lut_4_lut_LC_12_11_7  (
            .in0(N__36557),
            .in1(N__36449),
            .in2(N__36428),
            .in3(N__36319),
            .lcout(\Inst_core.Inst_controller.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Inst_core.Inst_controller.counter__i0_LC_12_12_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i0_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i0_LC_12_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i0_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__36275),
            .in2(_gnd_net_),
            .in3(N__36260),
            .lcout(\Inst_core.Inst_controller.counter_0 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\Inst_core.Inst_controller.n7845 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i1_LC_12_12_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i1_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i1_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i1_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__36257),
            .in2(_gnd_net_),
            .in3(N__36239),
            .lcout(\Inst_core.Inst_controller.counter_1 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7845 ),
            .carryout(\Inst_core.Inst_controller.n7846 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i2_LC_12_12_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i2_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i2_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i2_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__36236),
            .in2(_gnd_net_),
            .in3(N__36218),
            .lcout(\Inst_core.Inst_controller.counter_2 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7846 ),
            .carryout(\Inst_core.Inst_controller.n7847 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i3_LC_12_12_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i3_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i3_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i3_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__36204),
            .in2(_gnd_net_),
            .in3(N__36188),
            .lcout(\Inst_core.Inst_controller.counter_3 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7847 ),
            .carryout(\Inst_core.Inst_controller.n7848 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i4_LC_12_12_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i4_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i4_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i4_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__37100),
            .in2(_gnd_net_),
            .in3(N__37082),
            .lcout(\Inst_core.Inst_controller.counter_4 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7848 ),
            .carryout(\Inst_core.Inst_controller.n7849 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i5_LC_12_12_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i5_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i5_LC_12_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i5_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__37071),
            .in2(_gnd_net_),
            .in3(N__37055),
            .lcout(\Inst_core.Inst_controller.counter_5 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7849 ),
            .carryout(\Inst_core.Inst_controller.n7850 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i6_LC_12_12_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i6_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i6_LC_12_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i6_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__37044),
            .in2(_gnd_net_),
            .in3(N__37028),
            .lcout(\Inst_core.Inst_controller.counter_6 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7850 ),
            .carryout(\Inst_core.Inst_controller.n7851 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i7_LC_12_12_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i7_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i7_LC_12_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i7_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__37014),
            .in2(_gnd_net_),
            .in3(N__36992),
            .lcout(\Inst_core.Inst_controller.counter_7 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7851 ),
            .carryout(\Inst_core.Inst_controller.n7852 ),
            .clk(N__37612),
            .ce(N__37157),
            .sr(N__37116));
    defparam \Inst_core.Inst_controller.counter__i8_LC_12_13_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i8_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i8_LC_12_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i8_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__36978),
            .in2(_gnd_net_),
            .in3(N__36956),
            .lcout(\Inst_core.Inst_controller.counter_8 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\Inst_core.Inst_controller.n7853 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i9_LC_12_13_1 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i9_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i9_LC_12_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i9_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__36946),
            .in2(_gnd_net_),
            .in3(N__36932),
            .lcout(\Inst_core.Inst_controller.counter_9 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7853 ),
            .carryout(\Inst_core.Inst_controller.n7854 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i10_LC_12_13_2 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i10_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i10_LC_12_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i10_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__36921),
            .in2(_gnd_net_),
            .in3(N__36905),
            .lcout(\Inst_core.Inst_controller.counter_10 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7854 ),
            .carryout(\Inst_core.Inst_controller.n7855 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i11_LC_12_13_3 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i11_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i11_LC_12_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i11_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__36894),
            .in2(_gnd_net_),
            .in3(N__36878),
            .lcout(\Inst_core.Inst_controller.counter_11 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7855 ),
            .carryout(\Inst_core.Inst_controller.n7856 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i12_LC_12_13_4 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i12_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i12_LC_12_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i12_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__37789),
            .in2(_gnd_net_),
            .in3(N__37775),
            .lcout(\Inst_core.Inst_controller.counter_12 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7856 ),
            .carryout(\Inst_core.Inst_controller.n7857 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i13_LC_12_13_5 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i13_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i13_LC_12_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i13_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__37765),
            .in2(_gnd_net_),
            .in3(N__37751),
            .lcout(\Inst_core.Inst_controller.counter_13 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7857 ),
            .carryout(\Inst_core.Inst_controller.n7858 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i14_LC_12_13_6 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i14_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i14_LC_12_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i14_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__37741),
            .in2(_gnd_net_),
            .in3(N__37727),
            .lcout(\Inst_core.Inst_controller.counter_14 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7858 ),
            .carryout(\Inst_core.Inst_controller.n7859 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i15_LC_12_13_7 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i15_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i15_LC_12_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i15_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__37719),
            .in2(_gnd_net_),
            .in3(N__37700),
            .lcout(\Inst_core.Inst_controller.counter_15 ),
            .ltout(),
            .carryin(\Inst_core.Inst_controller.n7859 ),
            .carryout(\Inst_core.Inst_controller.n7860 ),
            .clk(N__37619),
            .ce(N__37156),
            .sr(N__37117));
    defparam \Inst_core.Inst_controller.counter__i16_LC_12_14_0 .C_ON=1'b1;
    defparam \Inst_core.Inst_controller.counter__i16_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i16_LC_12_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i16_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__37686),
            .in2(_gnd_net_),
            .in3(N__37670),
            .lcout(\Inst_core.Inst_controller.counter_16 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\Inst_core.Inst_controller.n7861 ),
            .clk(N__37625),
            .ce(N__37152),
            .sr(N__37124));
    defparam \Inst_core.Inst_controller.counter__i17_LC_12_14_1 .C_ON=1'b0;
    defparam \Inst_core.Inst_controller.counter__i17_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \Inst_core.Inst_controller.counter__i17_LC_12_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Inst_core.Inst_controller.counter__i17_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__37656),
            .in2(_gnd_net_),
            .in3(N__37667),
            .lcout(\Inst_core.Inst_controller.counter_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37625),
            .ce(N__37152),
            .sr(N__37124));
endmodule // la
